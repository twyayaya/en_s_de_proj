//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sat Jan 22 12:24:43 2022
// Version: v12.5 12.900.11.2
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// test1
module test1(
    // Inputs
    INn,
    clk,
    // Outputs
    ERRr,
    real_data
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  [71:0] INn;
input         clk;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output        ERRr;
output [63:0] real_data;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire          clk;
wire          ERRr_net_0;
wire   [71:0] INn;
wire   [63:0] real_data_net_0;
wire   [63:0] real_data_net_1;
wire          ERRr_net_1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign real_data_net_1 = real_data_net_0;
assign real_data[63:0] = real_data_net_1;
assign ERRr_net_1      = ERRr_net_0;
assign ERRr            = ERRr_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------de_v1
de_v1 de_v1_0(
        // Inputs
        .INn       ( INn ),
        .clk       ( clk ),
        // Outputs
        .ERRr      ( ERRr_net_0 ),
        .real_data ( real_data_net_0 ) 
        );


endmodule
