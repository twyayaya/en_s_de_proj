//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sat Jan 22 14:37:49 2022
// Version: v12.5 12.900.11.2
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// PF_TPSRAM_C0
module PF_TPSRAM_C0(
    // Inputs
    CLK,
    R_ADDR,
    R_EN,
    W_ADDR,
    W_DATA,
    W_EN,
    // Outputs
    R_DATA
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input         CLK;
input  [13:0] R_ADDR;
input         R_EN;
input  [13:0] W_ADDR;
input  [7:0]  W_DATA;
input         W_EN;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [7:0]  R_DATA;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire          CLK;
wire   [13:0] R_ADDR;
wire   [7:0]  R_DATA_0;
wire          R_EN;
wire   [13:0] W_ADDR;
wire   [7:0]  W_DATA;
wire          W_EN;
wire   [7:0]  R_DATA_0_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire          GND_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net    = 1'b0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign R_DATA_0_net_0 = R_DATA_0;
assign R_DATA[7:0]    = R_DATA_0_net_0;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM   -   Actel:SgCore:PF_TPSRAM:1.1.108
PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM PF_TPSRAM_C0_0(
        // Inputs
        .W_DATA ( W_DATA ),
        .W_ADDR ( W_ADDR ),
        .R_ADDR ( R_ADDR ),
        .W_EN   ( W_EN ),
        .R_EN   ( R_EN ),
        .CLK    ( CLK ),
        // Outputs
        .R_DATA ( R_DATA_0 ) 
        );


endmodule
