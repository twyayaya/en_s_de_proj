`timescale 1 ns/100 ps
// Version: v12.5 12.900.11.2


module PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM(
       W_DATA,
       R_DATA,
       W_ADDR,
       R_ADDR,
       W_EN,
       R_EN,
       CLK,
       WBYTE_EN
    );
input  [79:0] W_DATA;
output [79:0] R_DATA;
input  [13:0] W_ADDR;
input  [13:0] R_ADDR;
input  W_EN;
input  R_EN;
input  CLK;
input  [7:0] WBYTE_EN;

    wire \R_DATA_TEMPR0[0] , \R_DATA_TEMPR1[0] , \R_DATA_TEMPR2[0] , 
        \R_DATA_TEMPR3[0] , \R_DATA_TEMPR4[0] , \R_DATA_TEMPR5[0] , 
        \R_DATA_TEMPR6[0] , \R_DATA_TEMPR7[0] , \R_DATA_TEMPR8[0] , 
        \R_DATA_TEMPR9[0] , \R_DATA_TEMPR10[0] , \R_DATA_TEMPR11[0] , 
        \R_DATA_TEMPR12[0] , \R_DATA_TEMPR13[0] , \R_DATA_TEMPR14[0] , 
        \R_DATA_TEMPR15[0] , \R_DATA_TEMPR16[0] , \R_DATA_TEMPR17[0] , 
        \R_DATA_TEMPR18[0] , \R_DATA_TEMPR19[0] , \R_DATA_TEMPR20[0] , 
        \R_DATA_TEMPR21[0] , \R_DATA_TEMPR22[0] , \R_DATA_TEMPR23[0] , 
        \R_DATA_TEMPR24[0] , \R_DATA_TEMPR25[0] , \R_DATA_TEMPR26[0] , 
        \R_DATA_TEMPR27[0] , \R_DATA_TEMPR28[0] , \R_DATA_TEMPR29[0] , 
        \R_DATA_TEMPR30[0] , \R_DATA_TEMPR31[0] , \R_DATA_TEMPR0[1] , 
        \R_DATA_TEMPR1[1] , \R_DATA_TEMPR2[1] , \R_DATA_TEMPR3[1] , 
        \R_DATA_TEMPR4[1] , \R_DATA_TEMPR5[1] , \R_DATA_TEMPR6[1] , 
        \R_DATA_TEMPR7[1] , \R_DATA_TEMPR8[1] , \R_DATA_TEMPR9[1] , 
        \R_DATA_TEMPR10[1] , \R_DATA_TEMPR11[1] , \R_DATA_TEMPR12[1] , 
        \R_DATA_TEMPR13[1] , \R_DATA_TEMPR14[1] , \R_DATA_TEMPR15[1] , 
        \R_DATA_TEMPR16[1] , \R_DATA_TEMPR17[1] , \R_DATA_TEMPR18[1] , 
        \R_DATA_TEMPR19[1] , \R_DATA_TEMPR20[1] , \R_DATA_TEMPR21[1] , 
        \R_DATA_TEMPR22[1] , \R_DATA_TEMPR23[1] , \R_DATA_TEMPR24[1] , 
        \R_DATA_TEMPR25[1] , \R_DATA_TEMPR26[1] , \R_DATA_TEMPR27[1] , 
        \R_DATA_TEMPR28[1] , \R_DATA_TEMPR29[1] , \R_DATA_TEMPR30[1] , 
        \R_DATA_TEMPR31[1] , \R_DATA_TEMPR0[2] , \R_DATA_TEMPR1[2] , 
        \R_DATA_TEMPR2[2] , \R_DATA_TEMPR3[2] , \R_DATA_TEMPR4[2] , 
        \R_DATA_TEMPR5[2] , \R_DATA_TEMPR6[2] , \R_DATA_TEMPR7[2] , 
        \R_DATA_TEMPR8[2] , \R_DATA_TEMPR9[2] , \R_DATA_TEMPR10[2] , 
        \R_DATA_TEMPR11[2] , \R_DATA_TEMPR12[2] , \R_DATA_TEMPR13[2] , 
        \R_DATA_TEMPR14[2] , \R_DATA_TEMPR15[2] , \R_DATA_TEMPR16[2] , 
        \R_DATA_TEMPR17[2] , \R_DATA_TEMPR18[2] , \R_DATA_TEMPR19[2] , 
        \R_DATA_TEMPR20[2] , \R_DATA_TEMPR21[2] , \R_DATA_TEMPR22[2] , 
        \R_DATA_TEMPR23[2] , \R_DATA_TEMPR24[2] , \R_DATA_TEMPR25[2] , 
        \R_DATA_TEMPR26[2] , \R_DATA_TEMPR27[2] , \R_DATA_TEMPR28[2] , 
        \R_DATA_TEMPR29[2] , \R_DATA_TEMPR30[2] , \R_DATA_TEMPR31[2] , 
        \R_DATA_TEMPR0[3] , \R_DATA_TEMPR1[3] , \R_DATA_TEMPR2[3] , 
        \R_DATA_TEMPR3[3] , \R_DATA_TEMPR4[3] , \R_DATA_TEMPR5[3] , 
        \R_DATA_TEMPR6[3] , \R_DATA_TEMPR7[3] , \R_DATA_TEMPR8[3] , 
        \R_DATA_TEMPR9[3] , \R_DATA_TEMPR10[3] , \R_DATA_TEMPR11[3] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR13[3] , \R_DATA_TEMPR14[3] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR16[3] , \R_DATA_TEMPR17[3] , 
        \R_DATA_TEMPR18[3] , \R_DATA_TEMPR19[3] , \R_DATA_TEMPR20[3] , 
        \R_DATA_TEMPR21[3] , \R_DATA_TEMPR22[3] , \R_DATA_TEMPR23[3] , 
        \R_DATA_TEMPR24[3] , \R_DATA_TEMPR25[3] , \R_DATA_TEMPR26[3] , 
        \R_DATA_TEMPR27[3] , \R_DATA_TEMPR28[3] , \R_DATA_TEMPR29[3] , 
        \R_DATA_TEMPR30[3] , \R_DATA_TEMPR31[3] , \R_DATA_TEMPR0[4] , 
        \R_DATA_TEMPR1[4] , \R_DATA_TEMPR2[4] , \R_DATA_TEMPR3[4] , 
        \R_DATA_TEMPR4[4] , \R_DATA_TEMPR5[4] , \R_DATA_TEMPR6[4] , 
        \R_DATA_TEMPR7[4] , \R_DATA_TEMPR8[4] , \R_DATA_TEMPR9[4] , 
        \R_DATA_TEMPR10[4] , \R_DATA_TEMPR11[4] , \R_DATA_TEMPR12[4] , 
        \R_DATA_TEMPR13[4] , \R_DATA_TEMPR14[4] , \R_DATA_TEMPR15[4] , 
        \R_DATA_TEMPR16[4] , \R_DATA_TEMPR17[4] , \R_DATA_TEMPR18[4] , 
        \R_DATA_TEMPR19[4] , \R_DATA_TEMPR20[4] , \R_DATA_TEMPR21[4] , 
        \R_DATA_TEMPR22[4] , \R_DATA_TEMPR23[4] , \R_DATA_TEMPR24[4] , 
        \R_DATA_TEMPR25[4] , \R_DATA_TEMPR26[4] , \R_DATA_TEMPR27[4] , 
        \R_DATA_TEMPR28[4] , \R_DATA_TEMPR29[4] , \R_DATA_TEMPR30[4] , 
        \R_DATA_TEMPR31[4] , \R_DATA_TEMPR0[5] , \R_DATA_TEMPR1[5] , 
        \R_DATA_TEMPR2[5] , \R_DATA_TEMPR3[5] , \R_DATA_TEMPR4[5] , 
        \R_DATA_TEMPR5[5] , \R_DATA_TEMPR6[5] , \R_DATA_TEMPR7[5] , 
        \R_DATA_TEMPR8[5] , \R_DATA_TEMPR9[5] , \R_DATA_TEMPR10[5] , 
        \R_DATA_TEMPR11[5] , \R_DATA_TEMPR12[5] , \R_DATA_TEMPR13[5] , 
        \R_DATA_TEMPR14[5] , \R_DATA_TEMPR15[5] , \R_DATA_TEMPR16[5] , 
        \R_DATA_TEMPR17[5] , \R_DATA_TEMPR18[5] , \R_DATA_TEMPR19[5] , 
        \R_DATA_TEMPR20[5] , \R_DATA_TEMPR21[5] , \R_DATA_TEMPR22[5] , 
        \R_DATA_TEMPR23[5] , \R_DATA_TEMPR24[5] , \R_DATA_TEMPR25[5] , 
        \R_DATA_TEMPR26[5] , \R_DATA_TEMPR27[5] , \R_DATA_TEMPR28[5] , 
        \R_DATA_TEMPR29[5] , \R_DATA_TEMPR30[5] , \R_DATA_TEMPR31[5] , 
        \R_DATA_TEMPR0[6] , \R_DATA_TEMPR1[6] , \R_DATA_TEMPR2[6] , 
        \R_DATA_TEMPR3[6] , \R_DATA_TEMPR4[6] , \R_DATA_TEMPR5[6] , 
        \R_DATA_TEMPR6[6] , \R_DATA_TEMPR7[6] , \R_DATA_TEMPR8[6] , 
        \R_DATA_TEMPR9[6] , \R_DATA_TEMPR10[6] , \R_DATA_TEMPR11[6] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR13[6] , \R_DATA_TEMPR14[6] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR16[6] , \R_DATA_TEMPR17[6] , 
        \R_DATA_TEMPR18[6] , \R_DATA_TEMPR19[6] , \R_DATA_TEMPR20[6] , 
        \R_DATA_TEMPR21[6] , \R_DATA_TEMPR22[6] , \R_DATA_TEMPR23[6] , 
        \R_DATA_TEMPR24[6] , \R_DATA_TEMPR25[6] , \R_DATA_TEMPR26[6] , 
        \R_DATA_TEMPR27[6] , \R_DATA_TEMPR28[6] , \R_DATA_TEMPR29[6] , 
        \R_DATA_TEMPR30[6] , \R_DATA_TEMPR31[6] , \R_DATA_TEMPR0[7] , 
        \R_DATA_TEMPR1[7] , \R_DATA_TEMPR2[7] , \R_DATA_TEMPR3[7] , 
        \R_DATA_TEMPR4[7] , \R_DATA_TEMPR5[7] , \R_DATA_TEMPR6[7] , 
        \R_DATA_TEMPR7[7] , \R_DATA_TEMPR8[7] , \R_DATA_TEMPR9[7] , 
        \R_DATA_TEMPR10[7] , \R_DATA_TEMPR11[7] , \R_DATA_TEMPR12[7] , 
        \R_DATA_TEMPR13[7] , \R_DATA_TEMPR14[7] , \R_DATA_TEMPR15[7] , 
        \R_DATA_TEMPR16[7] , \R_DATA_TEMPR17[7] , \R_DATA_TEMPR18[7] , 
        \R_DATA_TEMPR19[7] , \R_DATA_TEMPR20[7] , \R_DATA_TEMPR21[7] , 
        \R_DATA_TEMPR22[7] , \R_DATA_TEMPR23[7] , \R_DATA_TEMPR24[7] , 
        \R_DATA_TEMPR25[7] , \R_DATA_TEMPR26[7] , \R_DATA_TEMPR27[7] , 
        \R_DATA_TEMPR28[7] , \R_DATA_TEMPR29[7] , \R_DATA_TEMPR30[7] , 
        \R_DATA_TEMPR31[7] , \R_DATA_TEMPR0[8] , \R_DATA_TEMPR1[8] , 
        \R_DATA_TEMPR2[8] , \R_DATA_TEMPR3[8] , \R_DATA_TEMPR4[8] , 
        \R_DATA_TEMPR5[8] , \R_DATA_TEMPR6[8] , \R_DATA_TEMPR7[8] , 
        \R_DATA_TEMPR8[8] , \R_DATA_TEMPR9[8] , \R_DATA_TEMPR10[8] , 
        \R_DATA_TEMPR11[8] , \R_DATA_TEMPR12[8] , \R_DATA_TEMPR13[8] , 
        \R_DATA_TEMPR14[8] , \R_DATA_TEMPR15[8] , \R_DATA_TEMPR16[8] , 
        \R_DATA_TEMPR17[8] , \R_DATA_TEMPR18[8] , \R_DATA_TEMPR19[8] , 
        \R_DATA_TEMPR20[8] , \R_DATA_TEMPR21[8] , \R_DATA_TEMPR22[8] , 
        \R_DATA_TEMPR23[8] , \R_DATA_TEMPR24[8] , \R_DATA_TEMPR25[8] , 
        \R_DATA_TEMPR26[8] , \R_DATA_TEMPR27[8] , \R_DATA_TEMPR28[8] , 
        \R_DATA_TEMPR29[8] , \R_DATA_TEMPR30[8] , \R_DATA_TEMPR31[8] , 
        \R_DATA_TEMPR0[9] , \R_DATA_TEMPR1[9] , \R_DATA_TEMPR2[9] , 
        \R_DATA_TEMPR3[9] , \R_DATA_TEMPR4[9] , \R_DATA_TEMPR5[9] , 
        \R_DATA_TEMPR6[9] , \R_DATA_TEMPR7[9] , \R_DATA_TEMPR8[9] , 
        \R_DATA_TEMPR9[9] , \R_DATA_TEMPR10[9] , \R_DATA_TEMPR11[9] , 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR13[9] , \R_DATA_TEMPR14[9] , 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR16[9] , \R_DATA_TEMPR17[9] , 
        \R_DATA_TEMPR18[9] , \R_DATA_TEMPR19[9] , \R_DATA_TEMPR20[9] , 
        \R_DATA_TEMPR21[9] , \R_DATA_TEMPR22[9] , \R_DATA_TEMPR23[9] , 
        \R_DATA_TEMPR24[9] , \R_DATA_TEMPR25[9] , \R_DATA_TEMPR26[9] , 
        \R_DATA_TEMPR27[9] , \R_DATA_TEMPR28[9] , \R_DATA_TEMPR29[9] , 
        \R_DATA_TEMPR30[9] , \R_DATA_TEMPR31[9] , \R_DATA_TEMPR0[10] , 
        \R_DATA_TEMPR1[10] , \R_DATA_TEMPR2[10] , \R_DATA_TEMPR3[10] , 
        \R_DATA_TEMPR4[10] , \R_DATA_TEMPR5[10] , \R_DATA_TEMPR6[10] , 
        \R_DATA_TEMPR7[10] , \R_DATA_TEMPR8[10] , \R_DATA_TEMPR9[10] , 
        \R_DATA_TEMPR10[10] , \R_DATA_TEMPR11[10] , 
        \R_DATA_TEMPR12[10] , \R_DATA_TEMPR13[10] , 
        \R_DATA_TEMPR14[10] , \R_DATA_TEMPR15[10] , 
        \R_DATA_TEMPR16[10] , \R_DATA_TEMPR17[10] , 
        \R_DATA_TEMPR18[10] , \R_DATA_TEMPR19[10] , 
        \R_DATA_TEMPR20[10] , \R_DATA_TEMPR21[10] , 
        \R_DATA_TEMPR22[10] , \R_DATA_TEMPR23[10] , 
        \R_DATA_TEMPR24[10] , \R_DATA_TEMPR25[10] , 
        \R_DATA_TEMPR26[10] , \R_DATA_TEMPR27[10] , 
        \R_DATA_TEMPR28[10] , \R_DATA_TEMPR29[10] , 
        \R_DATA_TEMPR30[10] , \R_DATA_TEMPR31[10] , 
        \R_DATA_TEMPR0[11] , \R_DATA_TEMPR1[11] , \R_DATA_TEMPR2[11] , 
        \R_DATA_TEMPR3[11] , \R_DATA_TEMPR4[11] , \R_DATA_TEMPR5[11] , 
        \R_DATA_TEMPR6[11] , \R_DATA_TEMPR7[11] , \R_DATA_TEMPR8[11] , 
        \R_DATA_TEMPR9[11] , \R_DATA_TEMPR10[11] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR12[11] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR14[11] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR16[11] , 
        \R_DATA_TEMPR17[11] , \R_DATA_TEMPR18[11] , 
        \R_DATA_TEMPR19[11] , \R_DATA_TEMPR20[11] , 
        \R_DATA_TEMPR21[11] , \R_DATA_TEMPR22[11] , 
        \R_DATA_TEMPR23[11] , \R_DATA_TEMPR24[11] , 
        \R_DATA_TEMPR25[11] , \R_DATA_TEMPR26[11] , 
        \R_DATA_TEMPR27[11] , \R_DATA_TEMPR28[11] , 
        \R_DATA_TEMPR29[11] , \R_DATA_TEMPR30[11] , 
        \R_DATA_TEMPR31[11] , \R_DATA_TEMPR0[12] , \R_DATA_TEMPR1[12] , 
        \R_DATA_TEMPR2[12] , \R_DATA_TEMPR3[12] , \R_DATA_TEMPR4[12] , 
        \R_DATA_TEMPR5[12] , \R_DATA_TEMPR6[12] , \R_DATA_TEMPR7[12] , 
        \R_DATA_TEMPR8[12] , \R_DATA_TEMPR9[12] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR11[12] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR13[12] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR15[12] , \R_DATA_TEMPR16[12] , 
        \R_DATA_TEMPR17[12] , \R_DATA_TEMPR18[12] , 
        \R_DATA_TEMPR19[12] , \R_DATA_TEMPR20[12] , 
        \R_DATA_TEMPR21[12] , \R_DATA_TEMPR22[12] , 
        \R_DATA_TEMPR23[12] , \R_DATA_TEMPR24[12] , 
        \R_DATA_TEMPR25[12] , \R_DATA_TEMPR26[12] , 
        \R_DATA_TEMPR27[12] , \R_DATA_TEMPR28[12] , 
        \R_DATA_TEMPR29[12] , \R_DATA_TEMPR30[12] , 
        \R_DATA_TEMPR31[12] , \R_DATA_TEMPR0[13] , \R_DATA_TEMPR1[13] , 
        \R_DATA_TEMPR2[13] , \R_DATA_TEMPR3[13] , \R_DATA_TEMPR4[13] , 
        \R_DATA_TEMPR5[13] , \R_DATA_TEMPR6[13] , \R_DATA_TEMPR7[13] , 
        \R_DATA_TEMPR8[13] , \R_DATA_TEMPR9[13] , \R_DATA_TEMPR10[13] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR12[13] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR14[13] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR16[13] , 
        \R_DATA_TEMPR17[13] , \R_DATA_TEMPR18[13] , 
        \R_DATA_TEMPR19[13] , \R_DATA_TEMPR20[13] , 
        \R_DATA_TEMPR21[13] , \R_DATA_TEMPR22[13] , 
        \R_DATA_TEMPR23[13] , \R_DATA_TEMPR24[13] , 
        \R_DATA_TEMPR25[13] , \R_DATA_TEMPR26[13] , 
        \R_DATA_TEMPR27[13] , \R_DATA_TEMPR28[13] , 
        \R_DATA_TEMPR29[13] , \R_DATA_TEMPR30[13] , 
        \R_DATA_TEMPR31[13] , \R_DATA_TEMPR0[14] , \R_DATA_TEMPR1[14] , 
        \R_DATA_TEMPR2[14] , \R_DATA_TEMPR3[14] , \R_DATA_TEMPR4[14] , 
        \R_DATA_TEMPR5[14] , \R_DATA_TEMPR6[14] , \R_DATA_TEMPR7[14] , 
        \R_DATA_TEMPR8[14] , \R_DATA_TEMPR9[14] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR11[14] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR13[14] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR15[14] , \R_DATA_TEMPR16[14] , 
        \R_DATA_TEMPR17[14] , \R_DATA_TEMPR18[14] , 
        \R_DATA_TEMPR19[14] , \R_DATA_TEMPR20[14] , 
        \R_DATA_TEMPR21[14] , \R_DATA_TEMPR22[14] , 
        \R_DATA_TEMPR23[14] , \R_DATA_TEMPR24[14] , 
        \R_DATA_TEMPR25[14] , \R_DATA_TEMPR26[14] , 
        \R_DATA_TEMPR27[14] , \R_DATA_TEMPR28[14] , 
        \R_DATA_TEMPR29[14] , \R_DATA_TEMPR30[14] , 
        \R_DATA_TEMPR31[14] , \R_DATA_TEMPR0[15] , \R_DATA_TEMPR1[15] , 
        \R_DATA_TEMPR2[15] , \R_DATA_TEMPR3[15] , \R_DATA_TEMPR4[15] , 
        \R_DATA_TEMPR5[15] , \R_DATA_TEMPR6[15] , \R_DATA_TEMPR7[15] , 
        \R_DATA_TEMPR8[15] , \R_DATA_TEMPR9[15] , \R_DATA_TEMPR10[15] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR12[15] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR14[15] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR16[15] , 
        \R_DATA_TEMPR17[15] , \R_DATA_TEMPR18[15] , 
        \R_DATA_TEMPR19[15] , \R_DATA_TEMPR20[15] , 
        \R_DATA_TEMPR21[15] , \R_DATA_TEMPR22[15] , 
        \R_DATA_TEMPR23[15] , \R_DATA_TEMPR24[15] , 
        \R_DATA_TEMPR25[15] , \R_DATA_TEMPR26[15] , 
        \R_DATA_TEMPR27[15] , \R_DATA_TEMPR28[15] , 
        \R_DATA_TEMPR29[15] , \R_DATA_TEMPR30[15] , 
        \R_DATA_TEMPR31[15] , \R_DATA_TEMPR0[16] , \R_DATA_TEMPR1[16] , 
        \R_DATA_TEMPR2[16] , \R_DATA_TEMPR3[16] , \R_DATA_TEMPR4[16] , 
        \R_DATA_TEMPR5[16] , \R_DATA_TEMPR6[16] , \R_DATA_TEMPR7[16] , 
        \R_DATA_TEMPR8[16] , \R_DATA_TEMPR9[16] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR11[16] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR13[16] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR15[16] , \R_DATA_TEMPR16[16] , 
        \R_DATA_TEMPR17[16] , \R_DATA_TEMPR18[16] , 
        \R_DATA_TEMPR19[16] , \R_DATA_TEMPR20[16] , 
        \R_DATA_TEMPR21[16] , \R_DATA_TEMPR22[16] , 
        \R_DATA_TEMPR23[16] , \R_DATA_TEMPR24[16] , 
        \R_DATA_TEMPR25[16] , \R_DATA_TEMPR26[16] , 
        \R_DATA_TEMPR27[16] , \R_DATA_TEMPR28[16] , 
        \R_DATA_TEMPR29[16] , \R_DATA_TEMPR30[16] , 
        \R_DATA_TEMPR31[16] , \R_DATA_TEMPR0[17] , \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR2[17] , \R_DATA_TEMPR3[17] , \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR5[17] , \R_DATA_TEMPR6[17] , \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR8[17] , \R_DATA_TEMPR9[17] , \R_DATA_TEMPR10[17] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR12[17] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR14[17] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR16[17] , 
        \R_DATA_TEMPR17[17] , \R_DATA_TEMPR18[17] , 
        \R_DATA_TEMPR19[17] , \R_DATA_TEMPR20[17] , 
        \R_DATA_TEMPR21[17] , \R_DATA_TEMPR22[17] , 
        \R_DATA_TEMPR23[17] , \R_DATA_TEMPR24[17] , 
        \R_DATA_TEMPR25[17] , \R_DATA_TEMPR26[17] , 
        \R_DATA_TEMPR27[17] , \R_DATA_TEMPR28[17] , 
        \R_DATA_TEMPR29[17] , \R_DATA_TEMPR30[17] , 
        \R_DATA_TEMPR31[17] , \R_DATA_TEMPR0[18] , \R_DATA_TEMPR1[18] , 
        \R_DATA_TEMPR2[18] , \R_DATA_TEMPR3[18] , \R_DATA_TEMPR4[18] , 
        \R_DATA_TEMPR5[18] , \R_DATA_TEMPR6[18] , \R_DATA_TEMPR7[18] , 
        \R_DATA_TEMPR8[18] , \R_DATA_TEMPR9[18] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR11[18] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR13[18] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR15[18] , \R_DATA_TEMPR16[18] , 
        \R_DATA_TEMPR17[18] , \R_DATA_TEMPR18[18] , 
        \R_DATA_TEMPR19[18] , \R_DATA_TEMPR20[18] , 
        \R_DATA_TEMPR21[18] , \R_DATA_TEMPR22[18] , 
        \R_DATA_TEMPR23[18] , \R_DATA_TEMPR24[18] , 
        \R_DATA_TEMPR25[18] , \R_DATA_TEMPR26[18] , 
        \R_DATA_TEMPR27[18] , \R_DATA_TEMPR28[18] , 
        \R_DATA_TEMPR29[18] , \R_DATA_TEMPR30[18] , 
        \R_DATA_TEMPR31[18] , \R_DATA_TEMPR0[19] , \R_DATA_TEMPR1[19] , 
        \R_DATA_TEMPR2[19] , \R_DATA_TEMPR3[19] , \R_DATA_TEMPR4[19] , 
        \R_DATA_TEMPR5[19] , \R_DATA_TEMPR6[19] , \R_DATA_TEMPR7[19] , 
        \R_DATA_TEMPR8[19] , \R_DATA_TEMPR9[19] , \R_DATA_TEMPR10[19] , 
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR12[19] , 
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR14[19] , 
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR16[19] , 
        \R_DATA_TEMPR17[19] , \R_DATA_TEMPR18[19] , 
        \R_DATA_TEMPR19[19] , \R_DATA_TEMPR20[19] , 
        \R_DATA_TEMPR21[19] , \R_DATA_TEMPR22[19] , 
        \R_DATA_TEMPR23[19] , \R_DATA_TEMPR24[19] , 
        \R_DATA_TEMPR25[19] , \R_DATA_TEMPR26[19] , 
        \R_DATA_TEMPR27[19] , \R_DATA_TEMPR28[19] , 
        \R_DATA_TEMPR29[19] , \R_DATA_TEMPR30[19] , 
        \R_DATA_TEMPR31[19] , \R_DATA_TEMPR0[20] , \R_DATA_TEMPR1[20] , 
        \R_DATA_TEMPR2[20] , \R_DATA_TEMPR3[20] , \R_DATA_TEMPR4[20] , 
        \R_DATA_TEMPR5[20] , \R_DATA_TEMPR6[20] , \R_DATA_TEMPR7[20] , 
        \R_DATA_TEMPR8[20] , \R_DATA_TEMPR9[20] , \R_DATA_TEMPR10[20] , 
        \R_DATA_TEMPR11[20] , \R_DATA_TEMPR12[20] , 
        \R_DATA_TEMPR13[20] , \R_DATA_TEMPR14[20] , 
        \R_DATA_TEMPR15[20] , \R_DATA_TEMPR16[20] , 
        \R_DATA_TEMPR17[20] , \R_DATA_TEMPR18[20] , 
        \R_DATA_TEMPR19[20] , \R_DATA_TEMPR20[20] , 
        \R_DATA_TEMPR21[20] , \R_DATA_TEMPR22[20] , 
        \R_DATA_TEMPR23[20] , \R_DATA_TEMPR24[20] , 
        \R_DATA_TEMPR25[20] , \R_DATA_TEMPR26[20] , 
        \R_DATA_TEMPR27[20] , \R_DATA_TEMPR28[20] , 
        \R_DATA_TEMPR29[20] , \R_DATA_TEMPR30[20] , 
        \R_DATA_TEMPR31[20] , \R_DATA_TEMPR0[21] , \R_DATA_TEMPR1[21] , 
        \R_DATA_TEMPR2[21] , \R_DATA_TEMPR3[21] , \R_DATA_TEMPR4[21] , 
        \R_DATA_TEMPR5[21] , \R_DATA_TEMPR6[21] , \R_DATA_TEMPR7[21] , 
        \R_DATA_TEMPR8[21] , \R_DATA_TEMPR9[21] , \R_DATA_TEMPR10[21] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR12[21] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR14[21] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR16[21] , 
        \R_DATA_TEMPR17[21] , \R_DATA_TEMPR18[21] , 
        \R_DATA_TEMPR19[21] , \R_DATA_TEMPR20[21] , 
        \R_DATA_TEMPR21[21] , \R_DATA_TEMPR22[21] , 
        \R_DATA_TEMPR23[21] , \R_DATA_TEMPR24[21] , 
        \R_DATA_TEMPR25[21] , \R_DATA_TEMPR26[21] , 
        \R_DATA_TEMPR27[21] , \R_DATA_TEMPR28[21] , 
        \R_DATA_TEMPR29[21] , \R_DATA_TEMPR30[21] , 
        \R_DATA_TEMPR31[21] , \R_DATA_TEMPR0[22] , \R_DATA_TEMPR1[22] , 
        \R_DATA_TEMPR2[22] , \R_DATA_TEMPR3[22] , \R_DATA_TEMPR4[22] , 
        \R_DATA_TEMPR5[22] , \R_DATA_TEMPR6[22] , \R_DATA_TEMPR7[22] , 
        \R_DATA_TEMPR8[22] , \R_DATA_TEMPR9[22] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR11[22] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR13[22] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR15[22] , \R_DATA_TEMPR16[22] , 
        \R_DATA_TEMPR17[22] , \R_DATA_TEMPR18[22] , 
        \R_DATA_TEMPR19[22] , \R_DATA_TEMPR20[22] , 
        \R_DATA_TEMPR21[22] , \R_DATA_TEMPR22[22] , 
        \R_DATA_TEMPR23[22] , \R_DATA_TEMPR24[22] , 
        \R_DATA_TEMPR25[22] , \R_DATA_TEMPR26[22] , 
        \R_DATA_TEMPR27[22] , \R_DATA_TEMPR28[22] , 
        \R_DATA_TEMPR29[22] , \R_DATA_TEMPR30[22] , 
        \R_DATA_TEMPR31[22] , \R_DATA_TEMPR0[23] , \R_DATA_TEMPR1[23] , 
        \R_DATA_TEMPR2[23] , \R_DATA_TEMPR3[23] , \R_DATA_TEMPR4[23] , 
        \R_DATA_TEMPR5[23] , \R_DATA_TEMPR6[23] , \R_DATA_TEMPR7[23] , 
        \R_DATA_TEMPR8[23] , \R_DATA_TEMPR9[23] , \R_DATA_TEMPR10[23] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR12[23] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR14[23] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR16[23] , 
        \R_DATA_TEMPR17[23] , \R_DATA_TEMPR18[23] , 
        \R_DATA_TEMPR19[23] , \R_DATA_TEMPR20[23] , 
        \R_DATA_TEMPR21[23] , \R_DATA_TEMPR22[23] , 
        \R_DATA_TEMPR23[23] , \R_DATA_TEMPR24[23] , 
        \R_DATA_TEMPR25[23] , \R_DATA_TEMPR26[23] , 
        \R_DATA_TEMPR27[23] , \R_DATA_TEMPR28[23] , 
        \R_DATA_TEMPR29[23] , \R_DATA_TEMPR30[23] , 
        \R_DATA_TEMPR31[23] , \R_DATA_TEMPR0[24] , \R_DATA_TEMPR1[24] , 
        \R_DATA_TEMPR2[24] , \R_DATA_TEMPR3[24] , \R_DATA_TEMPR4[24] , 
        \R_DATA_TEMPR5[24] , \R_DATA_TEMPR6[24] , \R_DATA_TEMPR7[24] , 
        \R_DATA_TEMPR8[24] , \R_DATA_TEMPR9[24] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR11[24] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR13[24] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR15[24] , \R_DATA_TEMPR16[24] , 
        \R_DATA_TEMPR17[24] , \R_DATA_TEMPR18[24] , 
        \R_DATA_TEMPR19[24] , \R_DATA_TEMPR20[24] , 
        \R_DATA_TEMPR21[24] , \R_DATA_TEMPR22[24] , 
        \R_DATA_TEMPR23[24] , \R_DATA_TEMPR24[24] , 
        \R_DATA_TEMPR25[24] , \R_DATA_TEMPR26[24] , 
        \R_DATA_TEMPR27[24] , \R_DATA_TEMPR28[24] , 
        \R_DATA_TEMPR29[24] , \R_DATA_TEMPR30[24] , 
        \R_DATA_TEMPR31[24] , \R_DATA_TEMPR0[25] , \R_DATA_TEMPR1[25] , 
        \R_DATA_TEMPR2[25] , \R_DATA_TEMPR3[25] , \R_DATA_TEMPR4[25] , 
        \R_DATA_TEMPR5[25] , \R_DATA_TEMPR6[25] , \R_DATA_TEMPR7[25] , 
        \R_DATA_TEMPR8[25] , \R_DATA_TEMPR9[25] , \R_DATA_TEMPR10[25] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR12[25] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR14[25] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR16[25] , 
        \R_DATA_TEMPR17[25] , \R_DATA_TEMPR18[25] , 
        \R_DATA_TEMPR19[25] , \R_DATA_TEMPR20[25] , 
        \R_DATA_TEMPR21[25] , \R_DATA_TEMPR22[25] , 
        \R_DATA_TEMPR23[25] , \R_DATA_TEMPR24[25] , 
        \R_DATA_TEMPR25[25] , \R_DATA_TEMPR26[25] , 
        \R_DATA_TEMPR27[25] , \R_DATA_TEMPR28[25] , 
        \R_DATA_TEMPR29[25] , \R_DATA_TEMPR30[25] , 
        \R_DATA_TEMPR31[25] , \R_DATA_TEMPR0[26] , \R_DATA_TEMPR1[26] , 
        \R_DATA_TEMPR2[26] , \R_DATA_TEMPR3[26] , \R_DATA_TEMPR4[26] , 
        \R_DATA_TEMPR5[26] , \R_DATA_TEMPR6[26] , \R_DATA_TEMPR7[26] , 
        \R_DATA_TEMPR8[26] , \R_DATA_TEMPR9[26] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR11[26] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR13[26] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR15[26] , \R_DATA_TEMPR16[26] , 
        \R_DATA_TEMPR17[26] , \R_DATA_TEMPR18[26] , 
        \R_DATA_TEMPR19[26] , \R_DATA_TEMPR20[26] , 
        \R_DATA_TEMPR21[26] , \R_DATA_TEMPR22[26] , 
        \R_DATA_TEMPR23[26] , \R_DATA_TEMPR24[26] , 
        \R_DATA_TEMPR25[26] , \R_DATA_TEMPR26[26] , 
        \R_DATA_TEMPR27[26] , \R_DATA_TEMPR28[26] , 
        \R_DATA_TEMPR29[26] , \R_DATA_TEMPR30[26] , 
        \R_DATA_TEMPR31[26] , \R_DATA_TEMPR0[27] , \R_DATA_TEMPR1[27] , 
        \R_DATA_TEMPR2[27] , \R_DATA_TEMPR3[27] , \R_DATA_TEMPR4[27] , 
        \R_DATA_TEMPR5[27] , \R_DATA_TEMPR6[27] , \R_DATA_TEMPR7[27] , 
        \R_DATA_TEMPR8[27] , \R_DATA_TEMPR9[27] , \R_DATA_TEMPR10[27] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR12[27] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR14[27] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR16[27] , 
        \R_DATA_TEMPR17[27] , \R_DATA_TEMPR18[27] , 
        \R_DATA_TEMPR19[27] , \R_DATA_TEMPR20[27] , 
        \R_DATA_TEMPR21[27] , \R_DATA_TEMPR22[27] , 
        \R_DATA_TEMPR23[27] , \R_DATA_TEMPR24[27] , 
        \R_DATA_TEMPR25[27] , \R_DATA_TEMPR26[27] , 
        \R_DATA_TEMPR27[27] , \R_DATA_TEMPR28[27] , 
        \R_DATA_TEMPR29[27] , \R_DATA_TEMPR30[27] , 
        \R_DATA_TEMPR31[27] , \R_DATA_TEMPR0[28] , \R_DATA_TEMPR1[28] , 
        \R_DATA_TEMPR2[28] , \R_DATA_TEMPR3[28] , \R_DATA_TEMPR4[28] , 
        \R_DATA_TEMPR5[28] , \R_DATA_TEMPR6[28] , \R_DATA_TEMPR7[28] , 
        \R_DATA_TEMPR8[28] , \R_DATA_TEMPR9[28] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR11[28] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR13[28] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR15[28] , \R_DATA_TEMPR16[28] , 
        \R_DATA_TEMPR17[28] , \R_DATA_TEMPR18[28] , 
        \R_DATA_TEMPR19[28] , \R_DATA_TEMPR20[28] , 
        \R_DATA_TEMPR21[28] , \R_DATA_TEMPR22[28] , 
        \R_DATA_TEMPR23[28] , \R_DATA_TEMPR24[28] , 
        \R_DATA_TEMPR25[28] , \R_DATA_TEMPR26[28] , 
        \R_DATA_TEMPR27[28] , \R_DATA_TEMPR28[28] , 
        \R_DATA_TEMPR29[28] , \R_DATA_TEMPR30[28] , 
        \R_DATA_TEMPR31[28] , \R_DATA_TEMPR0[29] , \R_DATA_TEMPR1[29] , 
        \R_DATA_TEMPR2[29] , \R_DATA_TEMPR3[29] , \R_DATA_TEMPR4[29] , 
        \R_DATA_TEMPR5[29] , \R_DATA_TEMPR6[29] , \R_DATA_TEMPR7[29] , 
        \R_DATA_TEMPR8[29] , \R_DATA_TEMPR9[29] , \R_DATA_TEMPR10[29] , 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR12[29] , 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR14[29] , 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR16[29] , 
        \R_DATA_TEMPR17[29] , \R_DATA_TEMPR18[29] , 
        \R_DATA_TEMPR19[29] , \R_DATA_TEMPR20[29] , 
        \R_DATA_TEMPR21[29] , \R_DATA_TEMPR22[29] , 
        \R_DATA_TEMPR23[29] , \R_DATA_TEMPR24[29] , 
        \R_DATA_TEMPR25[29] , \R_DATA_TEMPR26[29] , 
        \R_DATA_TEMPR27[29] , \R_DATA_TEMPR28[29] , 
        \R_DATA_TEMPR29[29] , \R_DATA_TEMPR30[29] , 
        \R_DATA_TEMPR31[29] , \R_DATA_TEMPR0[30] , \R_DATA_TEMPR1[30] , 
        \R_DATA_TEMPR2[30] , \R_DATA_TEMPR3[30] , \R_DATA_TEMPR4[30] , 
        \R_DATA_TEMPR5[30] , \R_DATA_TEMPR6[30] , \R_DATA_TEMPR7[30] , 
        \R_DATA_TEMPR8[30] , \R_DATA_TEMPR9[30] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR11[30] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR13[30] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR15[30] , \R_DATA_TEMPR16[30] , 
        \R_DATA_TEMPR17[30] , \R_DATA_TEMPR18[30] , 
        \R_DATA_TEMPR19[30] , \R_DATA_TEMPR20[30] , 
        \R_DATA_TEMPR21[30] , \R_DATA_TEMPR22[30] , 
        \R_DATA_TEMPR23[30] , \R_DATA_TEMPR24[30] , 
        \R_DATA_TEMPR25[30] , \R_DATA_TEMPR26[30] , 
        \R_DATA_TEMPR27[30] , \R_DATA_TEMPR28[30] , 
        \R_DATA_TEMPR29[30] , \R_DATA_TEMPR30[30] , 
        \R_DATA_TEMPR31[30] , \R_DATA_TEMPR0[31] , \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR2[31] , \R_DATA_TEMPR3[31] , \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR5[31] , \R_DATA_TEMPR6[31] , \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR8[31] , \R_DATA_TEMPR9[31] , \R_DATA_TEMPR10[31] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR12[31] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR14[31] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR16[31] , 
        \R_DATA_TEMPR17[31] , \R_DATA_TEMPR18[31] , 
        \R_DATA_TEMPR19[31] , \R_DATA_TEMPR20[31] , 
        \R_DATA_TEMPR21[31] , \R_DATA_TEMPR22[31] , 
        \R_DATA_TEMPR23[31] , \R_DATA_TEMPR24[31] , 
        \R_DATA_TEMPR25[31] , \R_DATA_TEMPR26[31] , 
        \R_DATA_TEMPR27[31] , \R_DATA_TEMPR28[31] , 
        \R_DATA_TEMPR29[31] , \R_DATA_TEMPR30[31] , 
        \R_DATA_TEMPR31[31] , \R_DATA_TEMPR0[32] , \R_DATA_TEMPR1[32] , 
        \R_DATA_TEMPR2[32] , \R_DATA_TEMPR3[32] , \R_DATA_TEMPR4[32] , 
        \R_DATA_TEMPR5[32] , \R_DATA_TEMPR6[32] , \R_DATA_TEMPR7[32] , 
        \R_DATA_TEMPR8[32] , \R_DATA_TEMPR9[32] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR11[32] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR13[32] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR15[32] , \R_DATA_TEMPR16[32] , 
        \R_DATA_TEMPR17[32] , \R_DATA_TEMPR18[32] , 
        \R_DATA_TEMPR19[32] , \R_DATA_TEMPR20[32] , 
        \R_DATA_TEMPR21[32] , \R_DATA_TEMPR22[32] , 
        \R_DATA_TEMPR23[32] , \R_DATA_TEMPR24[32] , 
        \R_DATA_TEMPR25[32] , \R_DATA_TEMPR26[32] , 
        \R_DATA_TEMPR27[32] , \R_DATA_TEMPR28[32] , 
        \R_DATA_TEMPR29[32] , \R_DATA_TEMPR30[32] , 
        \R_DATA_TEMPR31[32] , \R_DATA_TEMPR0[33] , \R_DATA_TEMPR1[33] , 
        \R_DATA_TEMPR2[33] , \R_DATA_TEMPR3[33] , \R_DATA_TEMPR4[33] , 
        \R_DATA_TEMPR5[33] , \R_DATA_TEMPR6[33] , \R_DATA_TEMPR7[33] , 
        \R_DATA_TEMPR8[33] , \R_DATA_TEMPR9[33] , \R_DATA_TEMPR10[33] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR12[33] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR14[33] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR16[33] , 
        \R_DATA_TEMPR17[33] , \R_DATA_TEMPR18[33] , 
        \R_DATA_TEMPR19[33] , \R_DATA_TEMPR20[33] , 
        \R_DATA_TEMPR21[33] , \R_DATA_TEMPR22[33] , 
        \R_DATA_TEMPR23[33] , \R_DATA_TEMPR24[33] , 
        \R_DATA_TEMPR25[33] , \R_DATA_TEMPR26[33] , 
        \R_DATA_TEMPR27[33] , \R_DATA_TEMPR28[33] , 
        \R_DATA_TEMPR29[33] , \R_DATA_TEMPR30[33] , 
        \R_DATA_TEMPR31[33] , \R_DATA_TEMPR0[34] , \R_DATA_TEMPR1[34] , 
        \R_DATA_TEMPR2[34] , \R_DATA_TEMPR3[34] , \R_DATA_TEMPR4[34] , 
        \R_DATA_TEMPR5[34] , \R_DATA_TEMPR6[34] , \R_DATA_TEMPR7[34] , 
        \R_DATA_TEMPR8[34] , \R_DATA_TEMPR9[34] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR11[34] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR13[34] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR15[34] , \R_DATA_TEMPR16[34] , 
        \R_DATA_TEMPR17[34] , \R_DATA_TEMPR18[34] , 
        \R_DATA_TEMPR19[34] , \R_DATA_TEMPR20[34] , 
        \R_DATA_TEMPR21[34] , \R_DATA_TEMPR22[34] , 
        \R_DATA_TEMPR23[34] , \R_DATA_TEMPR24[34] , 
        \R_DATA_TEMPR25[34] , \R_DATA_TEMPR26[34] , 
        \R_DATA_TEMPR27[34] , \R_DATA_TEMPR28[34] , 
        \R_DATA_TEMPR29[34] , \R_DATA_TEMPR30[34] , 
        \R_DATA_TEMPR31[34] , \R_DATA_TEMPR0[35] , \R_DATA_TEMPR1[35] , 
        \R_DATA_TEMPR2[35] , \R_DATA_TEMPR3[35] , \R_DATA_TEMPR4[35] , 
        \R_DATA_TEMPR5[35] , \R_DATA_TEMPR6[35] , \R_DATA_TEMPR7[35] , 
        \R_DATA_TEMPR8[35] , \R_DATA_TEMPR9[35] , \R_DATA_TEMPR10[35] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR12[35] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR14[35] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR16[35] , 
        \R_DATA_TEMPR17[35] , \R_DATA_TEMPR18[35] , 
        \R_DATA_TEMPR19[35] , \R_DATA_TEMPR20[35] , 
        \R_DATA_TEMPR21[35] , \R_DATA_TEMPR22[35] , 
        \R_DATA_TEMPR23[35] , \R_DATA_TEMPR24[35] , 
        \R_DATA_TEMPR25[35] , \R_DATA_TEMPR26[35] , 
        \R_DATA_TEMPR27[35] , \R_DATA_TEMPR28[35] , 
        \R_DATA_TEMPR29[35] , \R_DATA_TEMPR30[35] , 
        \R_DATA_TEMPR31[35] , \R_DATA_TEMPR0[36] , \R_DATA_TEMPR1[36] , 
        \R_DATA_TEMPR2[36] , \R_DATA_TEMPR3[36] , \R_DATA_TEMPR4[36] , 
        \R_DATA_TEMPR5[36] , \R_DATA_TEMPR6[36] , \R_DATA_TEMPR7[36] , 
        \R_DATA_TEMPR8[36] , \R_DATA_TEMPR9[36] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR11[36] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR13[36] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR15[36] , \R_DATA_TEMPR16[36] , 
        \R_DATA_TEMPR17[36] , \R_DATA_TEMPR18[36] , 
        \R_DATA_TEMPR19[36] , \R_DATA_TEMPR20[36] , 
        \R_DATA_TEMPR21[36] , \R_DATA_TEMPR22[36] , 
        \R_DATA_TEMPR23[36] , \R_DATA_TEMPR24[36] , 
        \R_DATA_TEMPR25[36] , \R_DATA_TEMPR26[36] , 
        \R_DATA_TEMPR27[36] , \R_DATA_TEMPR28[36] , 
        \R_DATA_TEMPR29[36] , \R_DATA_TEMPR30[36] , 
        \R_DATA_TEMPR31[36] , \R_DATA_TEMPR0[37] , \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR2[37] , \R_DATA_TEMPR3[37] , \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR5[37] , \R_DATA_TEMPR6[37] , \R_DATA_TEMPR7[37] , 
        \R_DATA_TEMPR8[37] , \R_DATA_TEMPR9[37] , \R_DATA_TEMPR10[37] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR12[37] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR14[37] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR16[37] , 
        \R_DATA_TEMPR17[37] , \R_DATA_TEMPR18[37] , 
        \R_DATA_TEMPR19[37] , \R_DATA_TEMPR20[37] , 
        \R_DATA_TEMPR21[37] , \R_DATA_TEMPR22[37] , 
        \R_DATA_TEMPR23[37] , \R_DATA_TEMPR24[37] , 
        \R_DATA_TEMPR25[37] , \R_DATA_TEMPR26[37] , 
        \R_DATA_TEMPR27[37] , \R_DATA_TEMPR28[37] , 
        \R_DATA_TEMPR29[37] , \R_DATA_TEMPR30[37] , 
        \R_DATA_TEMPR31[37] , \R_DATA_TEMPR0[38] , \R_DATA_TEMPR1[38] , 
        \R_DATA_TEMPR2[38] , \R_DATA_TEMPR3[38] , \R_DATA_TEMPR4[38] , 
        \R_DATA_TEMPR5[38] , \R_DATA_TEMPR6[38] , \R_DATA_TEMPR7[38] , 
        \R_DATA_TEMPR8[38] , \R_DATA_TEMPR9[38] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR11[38] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR13[38] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR15[38] , \R_DATA_TEMPR16[38] , 
        \R_DATA_TEMPR17[38] , \R_DATA_TEMPR18[38] , 
        \R_DATA_TEMPR19[38] , \R_DATA_TEMPR20[38] , 
        \R_DATA_TEMPR21[38] , \R_DATA_TEMPR22[38] , 
        \R_DATA_TEMPR23[38] , \R_DATA_TEMPR24[38] , 
        \R_DATA_TEMPR25[38] , \R_DATA_TEMPR26[38] , 
        \R_DATA_TEMPR27[38] , \R_DATA_TEMPR28[38] , 
        \R_DATA_TEMPR29[38] , \R_DATA_TEMPR30[38] , 
        \R_DATA_TEMPR31[38] , \R_DATA_TEMPR0[39] , \R_DATA_TEMPR1[39] , 
        \R_DATA_TEMPR2[39] , \R_DATA_TEMPR3[39] , \R_DATA_TEMPR4[39] , 
        \R_DATA_TEMPR5[39] , \R_DATA_TEMPR6[39] , \R_DATA_TEMPR7[39] , 
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR9[39] , \R_DATA_TEMPR10[39] , 
        \R_DATA_TEMPR11[39] , \R_DATA_TEMPR12[39] , 
        \R_DATA_TEMPR13[39] , \R_DATA_TEMPR14[39] , 
        \R_DATA_TEMPR15[39] , \R_DATA_TEMPR16[39] , 
        \R_DATA_TEMPR17[39] , \R_DATA_TEMPR18[39] , 
        \R_DATA_TEMPR19[39] , \R_DATA_TEMPR20[39] , 
        \R_DATA_TEMPR21[39] , \R_DATA_TEMPR22[39] , 
        \R_DATA_TEMPR23[39] , \R_DATA_TEMPR24[39] , 
        \R_DATA_TEMPR25[39] , \R_DATA_TEMPR26[39] , 
        \R_DATA_TEMPR27[39] , \R_DATA_TEMPR28[39] , 
        \R_DATA_TEMPR29[39] , \R_DATA_TEMPR30[39] , 
        \R_DATA_TEMPR31[39] , \R_DATA_TEMPR0[40] , \R_DATA_TEMPR1[40] , 
        \R_DATA_TEMPR2[40] , \R_DATA_TEMPR3[40] , \R_DATA_TEMPR4[40] , 
        \R_DATA_TEMPR5[40] , \R_DATA_TEMPR6[40] , \R_DATA_TEMPR7[40] , 
        \R_DATA_TEMPR8[40] , \R_DATA_TEMPR9[40] , \R_DATA_TEMPR10[40] , 
        \R_DATA_TEMPR11[40] , \R_DATA_TEMPR12[40] , 
        \R_DATA_TEMPR13[40] , \R_DATA_TEMPR14[40] , 
        \R_DATA_TEMPR15[40] , \R_DATA_TEMPR16[40] , 
        \R_DATA_TEMPR17[40] , \R_DATA_TEMPR18[40] , 
        \R_DATA_TEMPR19[40] , \R_DATA_TEMPR20[40] , 
        \R_DATA_TEMPR21[40] , \R_DATA_TEMPR22[40] , 
        \R_DATA_TEMPR23[40] , \R_DATA_TEMPR24[40] , 
        \R_DATA_TEMPR25[40] , \R_DATA_TEMPR26[40] , 
        \R_DATA_TEMPR27[40] , \R_DATA_TEMPR28[40] , 
        \R_DATA_TEMPR29[40] , \R_DATA_TEMPR30[40] , 
        \R_DATA_TEMPR31[40] , \R_DATA_TEMPR0[41] , \R_DATA_TEMPR1[41] , 
        \R_DATA_TEMPR2[41] , \R_DATA_TEMPR3[41] , \R_DATA_TEMPR4[41] , 
        \R_DATA_TEMPR5[41] , \R_DATA_TEMPR6[41] , \R_DATA_TEMPR7[41] , 
        \R_DATA_TEMPR8[41] , \R_DATA_TEMPR9[41] , \R_DATA_TEMPR10[41] , 
        \R_DATA_TEMPR11[41] , \R_DATA_TEMPR12[41] , 
        \R_DATA_TEMPR13[41] , \R_DATA_TEMPR14[41] , 
        \R_DATA_TEMPR15[41] , \R_DATA_TEMPR16[41] , 
        \R_DATA_TEMPR17[41] , \R_DATA_TEMPR18[41] , 
        \R_DATA_TEMPR19[41] , \R_DATA_TEMPR20[41] , 
        \R_DATA_TEMPR21[41] , \R_DATA_TEMPR22[41] , 
        \R_DATA_TEMPR23[41] , \R_DATA_TEMPR24[41] , 
        \R_DATA_TEMPR25[41] , \R_DATA_TEMPR26[41] , 
        \R_DATA_TEMPR27[41] , \R_DATA_TEMPR28[41] , 
        \R_DATA_TEMPR29[41] , \R_DATA_TEMPR30[41] , 
        \R_DATA_TEMPR31[41] , \R_DATA_TEMPR0[42] , \R_DATA_TEMPR1[42] , 
        \R_DATA_TEMPR2[42] , \R_DATA_TEMPR3[42] , \R_DATA_TEMPR4[42] , 
        \R_DATA_TEMPR5[42] , \R_DATA_TEMPR6[42] , \R_DATA_TEMPR7[42] , 
        \R_DATA_TEMPR8[42] , \R_DATA_TEMPR9[42] , \R_DATA_TEMPR10[42] , 
        \R_DATA_TEMPR11[42] , \R_DATA_TEMPR12[42] , 
        \R_DATA_TEMPR13[42] , \R_DATA_TEMPR14[42] , 
        \R_DATA_TEMPR15[42] , \R_DATA_TEMPR16[42] , 
        \R_DATA_TEMPR17[42] , \R_DATA_TEMPR18[42] , 
        \R_DATA_TEMPR19[42] , \R_DATA_TEMPR20[42] , 
        \R_DATA_TEMPR21[42] , \R_DATA_TEMPR22[42] , 
        \R_DATA_TEMPR23[42] , \R_DATA_TEMPR24[42] , 
        \R_DATA_TEMPR25[42] , \R_DATA_TEMPR26[42] , 
        \R_DATA_TEMPR27[42] , \R_DATA_TEMPR28[42] , 
        \R_DATA_TEMPR29[42] , \R_DATA_TEMPR30[42] , 
        \R_DATA_TEMPR31[42] , \R_DATA_TEMPR0[43] , \R_DATA_TEMPR1[43] , 
        \R_DATA_TEMPR2[43] , \R_DATA_TEMPR3[43] , \R_DATA_TEMPR4[43] , 
        \R_DATA_TEMPR5[43] , \R_DATA_TEMPR6[43] , \R_DATA_TEMPR7[43] , 
        \R_DATA_TEMPR8[43] , \R_DATA_TEMPR9[43] , \R_DATA_TEMPR10[43] , 
        \R_DATA_TEMPR11[43] , \R_DATA_TEMPR12[43] , 
        \R_DATA_TEMPR13[43] , \R_DATA_TEMPR14[43] , 
        \R_DATA_TEMPR15[43] , \R_DATA_TEMPR16[43] , 
        \R_DATA_TEMPR17[43] , \R_DATA_TEMPR18[43] , 
        \R_DATA_TEMPR19[43] , \R_DATA_TEMPR20[43] , 
        \R_DATA_TEMPR21[43] , \R_DATA_TEMPR22[43] , 
        \R_DATA_TEMPR23[43] , \R_DATA_TEMPR24[43] , 
        \R_DATA_TEMPR25[43] , \R_DATA_TEMPR26[43] , 
        \R_DATA_TEMPR27[43] , \R_DATA_TEMPR28[43] , 
        \R_DATA_TEMPR29[43] , \R_DATA_TEMPR30[43] , 
        \R_DATA_TEMPR31[43] , \R_DATA_TEMPR0[44] , \R_DATA_TEMPR1[44] , 
        \R_DATA_TEMPR2[44] , \R_DATA_TEMPR3[44] , \R_DATA_TEMPR4[44] , 
        \R_DATA_TEMPR5[44] , \R_DATA_TEMPR6[44] , \R_DATA_TEMPR7[44] , 
        \R_DATA_TEMPR8[44] , \R_DATA_TEMPR9[44] , \R_DATA_TEMPR10[44] , 
        \R_DATA_TEMPR11[44] , \R_DATA_TEMPR12[44] , 
        \R_DATA_TEMPR13[44] , \R_DATA_TEMPR14[44] , 
        \R_DATA_TEMPR15[44] , \R_DATA_TEMPR16[44] , 
        \R_DATA_TEMPR17[44] , \R_DATA_TEMPR18[44] , 
        \R_DATA_TEMPR19[44] , \R_DATA_TEMPR20[44] , 
        \R_DATA_TEMPR21[44] , \R_DATA_TEMPR22[44] , 
        \R_DATA_TEMPR23[44] , \R_DATA_TEMPR24[44] , 
        \R_DATA_TEMPR25[44] , \R_DATA_TEMPR26[44] , 
        \R_DATA_TEMPR27[44] , \R_DATA_TEMPR28[44] , 
        \R_DATA_TEMPR29[44] , \R_DATA_TEMPR30[44] , 
        \R_DATA_TEMPR31[44] , \R_DATA_TEMPR0[45] , \R_DATA_TEMPR1[45] , 
        \R_DATA_TEMPR2[45] , \R_DATA_TEMPR3[45] , \R_DATA_TEMPR4[45] , 
        \R_DATA_TEMPR5[45] , \R_DATA_TEMPR6[45] , \R_DATA_TEMPR7[45] , 
        \R_DATA_TEMPR8[45] , \R_DATA_TEMPR9[45] , \R_DATA_TEMPR10[45] , 
        \R_DATA_TEMPR11[45] , \R_DATA_TEMPR12[45] , 
        \R_DATA_TEMPR13[45] , \R_DATA_TEMPR14[45] , 
        \R_DATA_TEMPR15[45] , \R_DATA_TEMPR16[45] , 
        \R_DATA_TEMPR17[45] , \R_DATA_TEMPR18[45] , 
        \R_DATA_TEMPR19[45] , \R_DATA_TEMPR20[45] , 
        \R_DATA_TEMPR21[45] , \R_DATA_TEMPR22[45] , 
        \R_DATA_TEMPR23[45] , \R_DATA_TEMPR24[45] , 
        \R_DATA_TEMPR25[45] , \R_DATA_TEMPR26[45] , 
        \R_DATA_TEMPR27[45] , \R_DATA_TEMPR28[45] , 
        \R_DATA_TEMPR29[45] , \R_DATA_TEMPR30[45] , 
        \R_DATA_TEMPR31[45] , \R_DATA_TEMPR0[46] , \R_DATA_TEMPR1[46] , 
        \R_DATA_TEMPR2[46] , \R_DATA_TEMPR3[46] , \R_DATA_TEMPR4[46] , 
        \R_DATA_TEMPR5[46] , \R_DATA_TEMPR6[46] , \R_DATA_TEMPR7[46] , 
        \R_DATA_TEMPR8[46] , \R_DATA_TEMPR9[46] , \R_DATA_TEMPR10[46] , 
        \R_DATA_TEMPR11[46] , \R_DATA_TEMPR12[46] , 
        \R_DATA_TEMPR13[46] , \R_DATA_TEMPR14[46] , 
        \R_DATA_TEMPR15[46] , \R_DATA_TEMPR16[46] , 
        \R_DATA_TEMPR17[46] , \R_DATA_TEMPR18[46] , 
        \R_DATA_TEMPR19[46] , \R_DATA_TEMPR20[46] , 
        \R_DATA_TEMPR21[46] , \R_DATA_TEMPR22[46] , 
        \R_DATA_TEMPR23[46] , \R_DATA_TEMPR24[46] , 
        \R_DATA_TEMPR25[46] , \R_DATA_TEMPR26[46] , 
        \R_DATA_TEMPR27[46] , \R_DATA_TEMPR28[46] , 
        \R_DATA_TEMPR29[46] , \R_DATA_TEMPR30[46] , 
        \R_DATA_TEMPR31[46] , \R_DATA_TEMPR0[47] , \R_DATA_TEMPR1[47] , 
        \R_DATA_TEMPR2[47] , \R_DATA_TEMPR3[47] , \R_DATA_TEMPR4[47] , 
        \R_DATA_TEMPR5[47] , \R_DATA_TEMPR6[47] , \R_DATA_TEMPR7[47] , 
        \R_DATA_TEMPR8[47] , \R_DATA_TEMPR9[47] , \R_DATA_TEMPR10[47] , 
        \R_DATA_TEMPR11[47] , \R_DATA_TEMPR12[47] , 
        \R_DATA_TEMPR13[47] , \R_DATA_TEMPR14[47] , 
        \R_DATA_TEMPR15[47] , \R_DATA_TEMPR16[47] , 
        \R_DATA_TEMPR17[47] , \R_DATA_TEMPR18[47] , 
        \R_DATA_TEMPR19[47] , \R_DATA_TEMPR20[47] , 
        \R_DATA_TEMPR21[47] , \R_DATA_TEMPR22[47] , 
        \R_DATA_TEMPR23[47] , \R_DATA_TEMPR24[47] , 
        \R_DATA_TEMPR25[47] , \R_DATA_TEMPR26[47] , 
        \R_DATA_TEMPR27[47] , \R_DATA_TEMPR28[47] , 
        \R_DATA_TEMPR29[47] , \R_DATA_TEMPR30[47] , 
        \R_DATA_TEMPR31[47] , \R_DATA_TEMPR0[48] , \R_DATA_TEMPR1[48] , 
        \R_DATA_TEMPR2[48] , \R_DATA_TEMPR3[48] , \R_DATA_TEMPR4[48] , 
        \R_DATA_TEMPR5[48] , \R_DATA_TEMPR6[48] , \R_DATA_TEMPR7[48] , 
        \R_DATA_TEMPR8[48] , \R_DATA_TEMPR9[48] , \R_DATA_TEMPR10[48] , 
        \R_DATA_TEMPR11[48] , \R_DATA_TEMPR12[48] , 
        \R_DATA_TEMPR13[48] , \R_DATA_TEMPR14[48] , 
        \R_DATA_TEMPR15[48] , \R_DATA_TEMPR16[48] , 
        \R_DATA_TEMPR17[48] , \R_DATA_TEMPR18[48] , 
        \R_DATA_TEMPR19[48] , \R_DATA_TEMPR20[48] , 
        \R_DATA_TEMPR21[48] , \R_DATA_TEMPR22[48] , 
        \R_DATA_TEMPR23[48] , \R_DATA_TEMPR24[48] , 
        \R_DATA_TEMPR25[48] , \R_DATA_TEMPR26[48] , 
        \R_DATA_TEMPR27[48] , \R_DATA_TEMPR28[48] , 
        \R_DATA_TEMPR29[48] , \R_DATA_TEMPR30[48] , 
        \R_DATA_TEMPR31[48] , \R_DATA_TEMPR0[49] , \R_DATA_TEMPR1[49] , 
        \R_DATA_TEMPR2[49] , \R_DATA_TEMPR3[49] , \R_DATA_TEMPR4[49] , 
        \R_DATA_TEMPR5[49] , \R_DATA_TEMPR6[49] , \R_DATA_TEMPR7[49] , 
        \R_DATA_TEMPR8[49] , \R_DATA_TEMPR9[49] , \R_DATA_TEMPR10[49] , 
        \R_DATA_TEMPR11[49] , \R_DATA_TEMPR12[49] , 
        \R_DATA_TEMPR13[49] , \R_DATA_TEMPR14[49] , 
        \R_DATA_TEMPR15[49] , \R_DATA_TEMPR16[49] , 
        \R_DATA_TEMPR17[49] , \R_DATA_TEMPR18[49] , 
        \R_DATA_TEMPR19[49] , \R_DATA_TEMPR20[49] , 
        \R_DATA_TEMPR21[49] , \R_DATA_TEMPR22[49] , 
        \R_DATA_TEMPR23[49] , \R_DATA_TEMPR24[49] , 
        \R_DATA_TEMPR25[49] , \R_DATA_TEMPR26[49] , 
        \R_DATA_TEMPR27[49] , \R_DATA_TEMPR28[49] , 
        \R_DATA_TEMPR29[49] , \R_DATA_TEMPR30[49] , 
        \R_DATA_TEMPR31[49] , \R_DATA_TEMPR0[50] , \R_DATA_TEMPR1[50] , 
        \R_DATA_TEMPR2[50] , \R_DATA_TEMPR3[50] , \R_DATA_TEMPR4[50] , 
        \R_DATA_TEMPR5[50] , \R_DATA_TEMPR6[50] , \R_DATA_TEMPR7[50] , 
        \R_DATA_TEMPR8[50] , \R_DATA_TEMPR9[50] , \R_DATA_TEMPR10[50] , 
        \R_DATA_TEMPR11[50] , \R_DATA_TEMPR12[50] , 
        \R_DATA_TEMPR13[50] , \R_DATA_TEMPR14[50] , 
        \R_DATA_TEMPR15[50] , \R_DATA_TEMPR16[50] , 
        \R_DATA_TEMPR17[50] , \R_DATA_TEMPR18[50] , 
        \R_DATA_TEMPR19[50] , \R_DATA_TEMPR20[50] , 
        \R_DATA_TEMPR21[50] , \R_DATA_TEMPR22[50] , 
        \R_DATA_TEMPR23[50] , \R_DATA_TEMPR24[50] , 
        \R_DATA_TEMPR25[50] , \R_DATA_TEMPR26[50] , 
        \R_DATA_TEMPR27[50] , \R_DATA_TEMPR28[50] , 
        \R_DATA_TEMPR29[50] , \R_DATA_TEMPR30[50] , 
        \R_DATA_TEMPR31[50] , \R_DATA_TEMPR0[51] , \R_DATA_TEMPR1[51] , 
        \R_DATA_TEMPR2[51] , \R_DATA_TEMPR3[51] , \R_DATA_TEMPR4[51] , 
        \R_DATA_TEMPR5[51] , \R_DATA_TEMPR6[51] , \R_DATA_TEMPR7[51] , 
        \R_DATA_TEMPR8[51] , \R_DATA_TEMPR9[51] , \R_DATA_TEMPR10[51] , 
        \R_DATA_TEMPR11[51] , \R_DATA_TEMPR12[51] , 
        \R_DATA_TEMPR13[51] , \R_DATA_TEMPR14[51] , 
        \R_DATA_TEMPR15[51] , \R_DATA_TEMPR16[51] , 
        \R_DATA_TEMPR17[51] , \R_DATA_TEMPR18[51] , 
        \R_DATA_TEMPR19[51] , \R_DATA_TEMPR20[51] , 
        \R_DATA_TEMPR21[51] , \R_DATA_TEMPR22[51] , 
        \R_DATA_TEMPR23[51] , \R_DATA_TEMPR24[51] , 
        \R_DATA_TEMPR25[51] , \R_DATA_TEMPR26[51] , 
        \R_DATA_TEMPR27[51] , \R_DATA_TEMPR28[51] , 
        \R_DATA_TEMPR29[51] , \R_DATA_TEMPR30[51] , 
        \R_DATA_TEMPR31[51] , \R_DATA_TEMPR0[52] , \R_DATA_TEMPR1[52] , 
        \R_DATA_TEMPR2[52] , \R_DATA_TEMPR3[52] , \R_DATA_TEMPR4[52] , 
        \R_DATA_TEMPR5[52] , \R_DATA_TEMPR6[52] , \R_DATA_TEMPR7[52] , 
        \R_DATA_TEMPR8[52] , \R_DATA_TEMPR9[52] , \R_DATA_TEMPR10[52] , 
        \R_DATA_TEMPR11[52] , \R_DATA_TEMPR12[52] , 
        \R_DATA_TEMPR13[52] , \R_DATA_TEMPR14[52] , 
        \R_DATA_TEMPR15[52] , \R_DATA_TEMPR16[52] , 
        \R_DATA_TEMPR17[52] , \R_DATA_TEMPR18[52] , 
        \R_DATA_TEMPR19[52] , \R_DATA_TEMPR20[52] , 
        \R_DATA_TEMPR21[52] , \R_DATA_TEMPR22[52] , 
        \R_DATA_TEMPR23[52] , \R_DATA_TEMPR24[52] , 
        \R_DATA_TEMPR25[52] , \R_DATA_TEMPR26[52] , 
        \R_DATA_TEMPR27[52] , \R_DATA_TEMPR28[52] , 
        \R_DATA_TEMPR29[52] , \R_DATA_TEMPR30[52] , 
        \R_DATA_TEMPR31[52] , \R_DATA_TEMPR0[53] , \R_DATA_TEMPR1[53] , 
        \R_DATA_TEMPR2[53] , \R_DATA_TEMPR3[53] , \R_DATA_TEMPR4[53] , 
        \R_DATA_TEMPR5[53] , \R_DATA_TEMPR6[53] , \R_DATA_TEMPR7[53] , 
        \R_DATA_TEMPR8[53] , \R_DATA_TEMPR9[53] , \R_DATA_TEMPR10[53] , 
        \R_DATA_TEMPR11[53] , \R_DATA_TEMPR12[53] , 
        \R_DATA_TEMPR13[53] , \R_DATA_TEMPR14[53] , 
        \R_DATA_TEMPR15[53] , \R_DATA_TEMPR16[53] , 
        \R_DATA_TEMPR17[53] , \R_DATA_TEMPR18[53] , 
        \R_DATA_TEMPR19[53] , \R_DATA_TEMPR20[53] , 
        \R_DATA_TEMPR21[53] , \R_DATA_TEMPR22[53] , 
        \R_DATA_TEMPR23[53] , \R_DATA_TEMPR24[53] , 
        \R_DATA_TEMPR25[53] , \R_DATA_TEMPR26[53] , 
        \R_DATA_TEMPR27[53] , \R_DATA_TEMPR28[53] , 
        \R_DATA_TEMPR29[53] , \R_DATA_TEMPR30[53] , 
        \R_DATA_TEMPR31[53] , \R_DATA_TEMPR0[54] , \R_DATA_TEMPR1[54] , 
        \R_DATA_TEMPR2[54] , \R_DATA_TEMPR3[54] , \R_DATA_TEMPR4[54] , 
        \R_DATA_TEMPR5[54] , \R_DATA_TEMPR6[54] , \R_DATA_TEMPR7[54] , 
        \R_DATA_TEMPR8[54] , \R_DATA_TEMPR9[54] , \R_DATA_TEMPR10[54] , 
        \R_DATA_TEMPR11[54] , \R_DATA_TEMPR12[54] , 
        \R_DATA_TEMPR13[54] , \R_DATA_TEMPR14[54] , 
        \R_DATA_TEMPR15[54] , \R_DATA_TEMPR16[54] , 
        \R_DATA_TEMPR17[54] , \R_DATA_TEMPR18[54] , 
        \R_DATA_TEMPR19[54] , \R_DATA_TEMPR20[54] , 
        \R_DATA_TEMPR21[54] , \R_DATA_TEMPR22[54] , 
        \R_DATA_TEMPR23[54] , \R_DATA_TEMPR24[54] , 
        \R_DATA_TEMPR25[54] , \R_DATA_TEMPR26[54] , 
        \R_DATA_TEMPR27[54] , \R_DATA_TEMPR28[54] , 
        \R_DATA_TEMPR29[54] , \R_DATA_TEMPR30[54] , 
        \R_DATA_TEMPR31[54] , \R_DATA_TEMPR0[55] , \R_DATA_TEMPR1[55] , 
        \R_DATA_TEMPR2[55] , \R_DATA_TEMPR3[55] , \R_DATA_TEMPR4[55] , 
        \R_DATA_TEMPR5[55] , \R_DATA_TEMPR6[55] , \R_DATA_TEMPR7[55] , 
        \R_DATA_TEMPR8[55] , \R_DATA_TEMPR9[55] , \R_DATA_TEMPR10[55] , 
        \R_DATA_TEMPR11[55] , \R_DATA_TEMPR12[55] , 
        \R_DATA_TEMPR13[55] , \R_DATA_TEMPR14[55] , 
        \R_DATA_TEMPR15[55] , \R_DATA_TEMPR16[55] , 
        \R_DATA_TEMPR17[55] , \R_DATA_TEMPR18[55] , 
        \R_DATA_TEMPR19[55] , \R_DATA_TEMPR20[55] , 
        \R_DATA_TEMPR21[55] , \R_DATA_TEMPR22[55] , 
        \R_DATA_TEMPR23[55] , \R_DATA_TEMPR24[55] , 
        \R_DATA_TEMPR25[55] , \R_DATA_TEMPR26[55] , 
        \R_DATA_TEMPR27[55] , \R_DATA_TEMPR28[55] , 
        \R_DATA_TEMPR29[55] , \R_DATA_TEMPR30[55] , 
        \R_DATA_TEMPR31[55] , \R_DATA_TEMPR0[56] , \R_DATA_TEMPR1[56] , 
        \R_DATA_TEMPR2[56] , \R_DATA_TEMPR3[56] , \R_DATA_TEMPR4[56] , 
        \R_DATA_TEMPR5[56] , \R_DATA_TEMPR6[56] , \R_DATA_TEMPR7[56] , 
        \R_DATA_TEMPR8[56] , \R_DATA_TEMPR9[56] , \R_DATA_TEMPR10[56] , 
        \R_DATA_TEMPR11[56] , \R_DATA_TEMPR12[56] , 
        \R_DATA_TEMPR13[56] , \R_DATA_TEMPR14[56] , 
        \R_DATA_TEMPR15[56] , \R_DATA_TEMPR16[56] , 
        \R_DATA_TEMPR17[56] , \R_DATA_TEMPR18[56] , 
        \R_DATA_TEMPR19[56] , \R_DATA_TEMPR20[56] , 
        \R_DATA_TEMPR21[56] , \R_DATA_TEMPR22[56] , 
        \R_DATA_TEMPR23[56] , \R_DATA_TEMPR24[56] , 
        \R_DATA_TEMPR25[56] , \R_DATA_TEMPR26[56] , 
        \R_DATA_TEMPR27[56] , \R_DATA_TEMPR28[56] , 
        \R_DATA_TEMPR29[56] , \R_DATA_TEMPR30[56] , 
        \R_DATA_TEMPR31[56] , \R_DATA_TEMPR0[57] , \R_DATA_TEMPR1[57] , 
        \R_DATA_TEMPR2[57] , \R_DATA_TEMPR3[57] , \R_DATA_TEMPR4[57] , 
        \R_DATA_TEMPR5[57] , \R_DATA_TEMPR6[57] , \R_DATA_TEMPR7[57] , 
        \R_DATA_TEMPR8[57] , \R_DATA_TEMPR9[57] , \R_DATA_TEMPR10[57] , 
        \R_DATA_TEMPR11[57] , \R_DATA_TEMPR12[57] , 
        \R_DATA_TEMPR13[57] , \R_DATA_TEMPR14[57] , 
        \R_DATA_TEMPR15[57] , \R_DATA_TEMPR16[57] , 
        \R_DATA_TEMPR17[57] , \R_DATA_TEMPR18[57] , 
        \R_DATA_TEMPR19[57] , \R_DATA_TEMPR20[57] , 
        \R_DATA_TEMPR21[57] , \R_DATA_TEMPR22[57] , 
        \R_DATA_TEMPR23[57] , \R_DATA_TEMPR24[57] , 
        \R_DATA_TEMPR25[57] , \R_DATA_TEMPR26[57] , 
        \R_DATA_TEMPR27[57] , \R_DATA_TEMPR28[57] , 
        \R_DATA_TEMPR29[57] , \R_DATA_TEMPR30[57] , 
        \R_DATA_TEMPR31[57] , \R_DATA_TEMPR0[58] , \R_DATA_TEMPR1[58] , 
        \R_DATA_TEMPR2[58] , \R_DATA_TEMPR3[58] , \R_DATA_TEMPR4[58] , 
        \R_DATA_TEMPR5[58] , \R_DATA_TEMPR6[58] , \R_DATA_TEMPR7[58] , 
        \R_DATA_TEMPR8[58] , \R_DATA_TEMPR9[58] , \R_DATA_TEMPR10[58] , 
        \R_DATA_TEMPR11[58] , \R_DATA_TEMPR12[58] , 
        \R_DATA_TEMPR13[58] , \R_DATA_TEMPR14[58] , 
        \R_DATA_TEMPR15[58] , \R_DATA_TEMPR16[58] , 
        \R_DATA_TEMPR17[58] , \R_DATA_TEMPR18[58] , 
        \R_DATA_TEMPR19[58] , \R_DATA_TEMPR20[58] , 
        \R_DATA_TEMPR21[58] , \R_DATA_TEMPR22[58] , 
        \R_DATA_TEMPR23[58] , \R_DATA_TEMPR24[58] , 
        \R_DATA_TEMPR25[58] , \R_DATA_TEMPR26[58] , 
        \R_DATA_TEMPR27[58] , \R_DATA_TEMPR28[58] , 
        \R_DATA_TEMPR29[58] , \R_DATA_TEMPR30[58] , 
        \R_DATA_TEMPR31[58] , \R_DATA_TEMPR0[59] , \R_DATA_TEMPR1[59] , 
        \R_DATA_TEMPR2[59] , \R_DATA_TEMPR3[59] , \R_DATA_TEMPR4[59] , 
        \R_DATA_TEMPR5[59] , \R_DATA_TEMPR6[59] , \R_DATA_TEMPR7[59] , 
        \R_DATA_TEMPR8[59] , \R_DATA_TEMPR9[59] , \R_DATA_TEMPR10[59] , 
        \R_DATA_TEMPR11[59] , \R_DATA_TEMPR12[59] , 
        \R_DATA_TEMPR13[59] , \R_DATA_TEMPR14[59] , 
        \R_DATA_TEMPR15[59] , \R_DATA_TEMPR16[59] , 
        \R_DATA_TEMPR17[59] , \R_DATA_TEMPR18[59] , 
        \R_DATA_TEMPR19[59] , \R_DATA_TEMPR20[59] , 
        \R_DATA_TEMPR21[59] , \R_DATA_TEMPR22[59] , 
        \R_DATA_TEMPR23[59] , \R_DATA_TEMPR24[59] , 
        \R_DATA_TEMPR25[59] , \R_DATA_TEMPR26[59] , 
        \R_DATA_TEMPR27[59] , \R_DATA_TEMPR28[59] , 
        \R_DATA_TEMPR29[59] , \R_DATA_TEMPR30[59] , 
        \R_DATA_TEMPR31[59] , \R_DATA_TEMPR0[60] , \R_DATA_TEMPR1[60] , 
        \R_DATA_TEMPR2[60] , \R_DATA_TEMPR3[60] , \R_DATA_TEMPR4[60] , 
        \R_DATA_TEMPR5[60] , \R_DATA_TEMPR6[60] , \R_DATA_TEMPR7[60] , 
        \R_DATA_TEMPR8[60] , \R_DATA_TEMPR9[60] , \R_DATA_TEMPR10[60] , 
        \R_DATA_TEMPR11[60] , \R_DATA_TEMPR12[60] , 
        \R_DATA_TEMPR13[60] , \R_DATA_TEMPR14[60] , 
        \R_DATA_TEMPR15[60] , \R_DATA_TEMPR16[60] , 
        \R_DATA_TEMPR17[60] , \R_DATA_TEMPR18[60] , 
        \R_DATA_TEMPR19[60] , \R_DATA_TEMPR20[60] , 
        \R_DATA_TEMPR21[60] , \R_DATA_TEMPR22[60] , 
        \R_DATA_TEMPR23[60] , \R_DATA_TEMPR24[60] , 
        \R_DATA_TEMPR25[60] , \R_DATA_TEMPR26[60] , 
        \R_DATA_TEMPR27[60] , \R_DATA_TEMPR28[60] , 
        \R_DATA_TEMPR29[60] , \R_DATA_TEMPR30[60] , 
        \R_DATA_TEMPR31[60] , \R_DATA_TEMPR0[61] , \R_DATA_TEMPR1[61] , 
        \R_DATA_TEMPR2[61] , \R_DATA_TEMPR3[61] , \R_DATA_TEMPR4[61] , 
        \R_DATA_TEMPR5[61] , \R_DATA_TEMPR6[61] , \R_DATA_TEMPR7[61] , 
        \R_DATA_TEMPR8[61] , \R_DATA_TEMPR9[61] , \R_DATA_TEMPR10[61] , 
        \R_DATA_TEMPR11[61] , \R_DATA_TEMPR12[61] , 
        \R_DATA_TEMPR13[61] , \R_DATA_TEMPR14[61] , 
        \R_DATA_TEMPR15[61] , \R_DATA_TEMPR16[61] , 
        \R_DATA_TEMPR17[61] , \R_DATA_TEMPR18[61] , 
        \R_DATA_TEMPR19[61] , \R_DATA_TEMPR20[61] , 
        \R_DATA_TEMPR21[61] , \R_DATA_TEMPR22[61] , 
        \R_DATA_TEMPR23[61] , \R_DATA_TEMPR24[61] , 
        \R_DATA_TEMPR25[61] , \R_DATA_TEMPR26[61] , 
        \R_DATA_TEMPR27[61] , \R_DATA_TEMPR28[61] , 
        \R_DATA_TEMPR29[61] , \R_DATA_TEMPR30[61] , 
        \R_DATA_TEMPR31[61] , \R_DATA_TEMPR0[62] , \R_DATA_TEMPR1[62] , 
        \R_DATA_TEMPR2[62] , \R_DATA_TEMPR3[62] , \R_DATA_TEMPR4[62] , 
        \R_DATA_TEMPR5[62] , \R_DATA_TEMPR6[62] , \R_DATA_TEMPR7[62] , 
        \R_DATA_TEMPR8[62] , \R_DATA_TEMPR9[62] , \R_DATA_TEMPR10[62] , 
        \R_DATA_TEMPR11[62] , \R_DATA_TEMPR12[62] , 
        \R_DATA_TEMPR13[62] , \R_DATA_TEMPR14[62] , 
        \R_DATA_TEMPR15[62] , \R_DATA_TEMPR16[62] , 
        \R_DATA_TEMPR17[62] , \R_DATA_TEMPR18[62] , 
        \R_DATA_TEMPR19[62] , \R_DATA_TEMPR20[62] , 
        \R_DATA_TEMPR21[62] , \R_DATA_TEMPR22[62] , 
        \R_DATA_TEMPR23[62] , \R_DATA_TEMPR24[62] , 
        \R_DATA_TEMPR25[62] , \R_DATA_TEMPR26[62] , 
        \R_DATA_TEMPR27[62] , \R_DATA_TEMPR28[62] , 
        \R_DATA_TEMPR29[62] , \R_DATA_TEMPR30[62] , 
        \R_DATA_TEMPR31[62] , \R_DATA_TEMPR0[63] , \R_DATA_TEMPR1[63] , 
        \R_DATA_TEMPR2[63] , \R_DATA_TEMPR3[63] , \R_DATA_TEMPR4[63] , 
        \R_DATA_TEMPR5[63] , \R_DATA_TEMPR6[63] , \R_DATA_TEMPR7[63] , 
        \R_DATA_TEMPR8[63] , \R_DATA_TEMPR9[63] , \R_DATA_TEMPR10[63] , 
        \R_DATA_TEMPR11[63] , \R_DATA_TEMPR12[63] , 
        \R_DATA_TEMPR13[63] , \R_DATA_TEMPR14[63] , 
        \R_DATA_TEMPR15[63] , \R_DATA_TEMPR16[63] , 
        \R_DATA_TEMPR17[63] , \R_DATA_TEMPR18[63] , 
        \R_DATA_TEMPR19[63] , \R_DATA_TEMPR20[63] , 
        \R_DATA_TEMPR21[63] , \R_DATA_TEMPR22[63] , 
        \R_DATA_TEMPR23[63] , \R_DATA_TEMPR24[63] , 
        \R_DATA_TEMPR25[63] , \R_DATA_TEMPR26[63] , 
        \R_DATA_TEMPR27[63] , \R_DATA_TEMPR28[63] , 
        \R_DATA_TEMPR29[63] , \R_DATA_TEMPR30[63] , 
        \R_DATA_TEMPR31[63] , \R_DATA_TEMPR0[64] , \R_DATA_TEMPR1[64] , 
        \R_DATA_TEMPR2[64] , \R_DATA_TEMPR3[64] , \R_DATA_TEMPR4[64] , 
        \R_DATA_TEMPR5[64] , \R_DATA_TEMPR6[64] , \R_DATA_TEMPR7[64] , 
        \R_DATA_TEMPR8[64] , \R_DATA_TEMPR9[64] , \R_DATA_TEMPR10[64] , 
        \R_DATA_TEMPR11[64] , \R_DATA_TEMPR12[64] , 
        \R_DATA_TEMPR13[64] , \R_DATA_TEMPR14[64] , 
        \R_DATA_TEMPR15[64] , \R_DATA_TEMPR16[64] , 
        \R_DATA_TEMPR17[64] , \R_DATA_TEMPR18[64] , 
        \R_DATA_TEMPR19[64] , \R_DATA_TEMPR20[64] , 
        \R_DATA_TEMPR21[64] , \R_DATA_TEMPR22[64] , 
        \R_DATA_TEMPR23[64] , \R_DATA_TEMPR24[64] , 
        \R_DATA_TEMPR25[64] , \R_DATA_TEMPR26[64] , 
        \R_DATA_TEMPR27[64] , \R_DATA_TEMPR28[64] , 
        \R_DATA_TEMPR29[64] , \R_DATA_TEMPR30[64] , 
        \R_DATA_TEMPR31[64] , \R_DATA_TEMPR0[65] , \R_DATA_TEMPR1[65] , 
        \R_DATA_TEMPR2[65] , \R_DATA_TEMPR3[65] , \R_DATA_TEMPR4[65] , 
        \R_DATA_TEMPR5[65] , \R_DATA_TEMPR6[65] , \R_DATA_TEMPR7[65] , 
        \R_DATA_TEMPR8[65] , \R_DATA_TEMPR9[65] , \R_DATA_TEMPR10[65] , 
        \R_DATA_TEMPR11[65] , \R_DATA_TEMPR12[65] , 
        \R_DATA_TEMPR13[65] , \R_DATA_TEMPR14[65] , 
        \R_DATA_TEMPR15[65] , \R_DATA_TEMPR16[65] , 
        \R_DATA_TEMPR17[65] , \R_DATA_TEMPR18[65] , 
        \R_DATA_TEMPR19[65] , \R_DATA_TEMPR20[65] , 
        \R_DATA_TEMPR21[65] , \R_DATA_TEMPR22[65] , 
        \R_DATA_TEMPR23[65] , \R_DATA_TEMPR24[65] , 
        \R_DATA_TEMPR25[65] , \R_DATA_TEMPR26[65] , 
        \R_DATA_TEMPR27[65] , \R_DATA_TEMPR28[65] , 
        \R_DATA_TEMPR29[65] , \R_DATA_TEMPR30[65] , 
        \R_DATA_TEMPR31[65] , \R_DATA_TEMPR0[66] , \R_DATA_TEMPR1[66] , 
        \R_DATA_TEMPR2[66] , \R_DATA_TEMPR3[66] , \R_DATA_TEMPR4[66] , 
        \R_DATA_TEMPR5[66] , \R_DATA_TEMPR6[66] , \R_DATA_TEMPR7[66] , 
        \R_DATA_TEMPR8[66] , \R_DATA_TEMPR9[66] , \R_DATA_TEMPR10[66] , 
        \R_DATA_TEMPR11[66] , \R_DATA_TEMPR12[66] , 
        \R_DATA_TEMPR13[66] , \R_DATA_TEMPR14[66] , 
        \R_DATA_TEMPR15[66] , \R_DATA_TEMPR16[66] , 
        \R_DATA_TEMPR17[66] , \R_DATA_TEMPR18[66] , 
        \R_DATA_TEMPR19[66] , \R_DATA_TEMPR20[66] , 
        \R_DATA_TEMPR21[66] , \R_DATA_TEMPR22[66] , 
        \R_DATA_TEMPR23[66] , \R_DATA_TEMPR24[66] , 
        \R_DATA_TEMPR25[66] , \R_DATA_TEMPR26[66] , 
        \R_DATA_TEMPR27[66] , \R_DATA_TEMPR28[66] , 
        \R_DATA_TEMPR29[66] , \R_DATA_TEMPR30[66] , 
        \R_DATA_TEMPR31[66] , \R_DATA_TEMPR0[67] , \R_DATA_TEMPR1[67] , 
        \R_DATA_TEMPR2[67] , \R_DATA_TEMPR3[67] , \R_DATA_TEMPR4[67] , 
        \R_DATA_TEMPR5[67] , \R_DATA_TEMPR6[67] , \R_DATA_TEMPR7[67] , 
        \R_DATA_TEMPR8[67] , \R_DATA_TEMPR9[67] , \R_DATA_TEMPR10[67] , 
        \R_DATA_TEMPR11[67] , \R_DATA_TEMPR12[67] , 
        \R_DATA_TEMPR13[67] , \R_DATA_TEMPR14[67] , 
        \R_DATA_TEMPR15[67] , \R_DATA_TEMPR16[67] , 
        \R_DATA_TEMPR17[67] , \R_DATA_TEMPR18[67] , 
        \R_DATA_TEMPR19[67] , \R_DATA_TEMPR20[67] , 
        \R_DATA_TEMPR21[67] , \R_DATA_TEMPR22[67] , 
        \R_DATA_TEMPR23[67] , \R_DATA_TEMPR24[67] , 
        \R_DATA_TEMPR25[67] , \R_DATA_TEMPR26[67] , 
        \R_DATA_TEMPR27[67] , \R_DATA_TEMPR28[67] , 
        \R_DATA_TEMPR29[67] , \R_DATA_TEMPR30[67] , 
        \R_DATA_TEMPR31[67] , \R_DATA_TEMPR0[68] , \R_DATA_TEMPR1[68] , 
        \R_DATA_TEMPR2[68] , \R_DATA_TEMPR3[68] , \R_DATA_TEMPR4[68] , 
        \R_DATA_TEMPR5[68] , \R_DATA_TEMPR6[68] , \R_DATA_TEMPR7[68] , 
        \R_DATA_TEMPR8[68] , \R_DATA_TEMPR9[68] , \R_DATA_TEMPR10[68] , 
        \R_DATA_TEMPR11[68] , \R_DATA_TEMPR12[68] , 
        \R_DATA_TEMPR13[68] , \R_DATA_TEMPR14[68] , 
        \R_DATA_TEMPR15[68] , \R_DATA_TEMPR16[68] , 
        \R_DATA_TEMPR17[68] , \R_DATA_TEMPR18[68] , 
        \R_DATA_TEMPR19[68] , \R_DATA_TEMPR20[68] , 
        \R_DATA_TEMPR21[68] , \R_DATA_TEMPR22[68] , 
        \R_DATA_TEMPR23[68] , \R_DATA_TEMPR24[68] , 
        \R_DATA_TEMPR25[68] , \R_DATA_TEMPR26[68] , 
        \R_DATA_TEMPR27[68] , \R_DATA_TEMPR28[68] , 
        \R_DATA_TEMPR29[68] , \R_DATA_TEMPR30[68] , 
        \R_DATA_TEMPR31[68] , \R_DATA_TEMPR0[69] , \R_DATA_TEMPR1[69] , 
        \R_DATA_TEMPR2[69] , \R_DATA_TEMPR3[69] , \R_DATA_TEMPR4[69] , 
        \R_DATA_TEMPR5[69] , \R_DATA_TEMPR6[69] , \R_DATA_TEMPR7[69] , 
        \R_DATA_TEMPR8[69] , \R_DATA_TEMPR9[69] , \R_DATA_TEMPR10[69] , 
        \R_DATA_TEMPR11[69] , \R_DATA_TEMPR12[69] , 
        \R_DATA_TEMPR13[69] , \R_DATA_TEMPR14[69] , 
        \R_DATA_TEMPR15[69] , \R_DATA_TEMPR16[69] , 
        \R_DATA_TEMPR17[69] , \R_DATA_TEMPR18[69] , 
        \R_DATA_TEMPR19[69] , \R_DATA_TEMPR20[69] , 
        \R_DATA_TEMPR21[69] , \R_DATA_TEMPR22[69] , 
        \R_DATA_TEMPR23[69] , \R_DATA_TEMPR24[69] , 
        \R_DATA_TEMPR25[69] , \R_DATA_TEMPR26[69] , 
        \R_DATA_TEMPR27[69] , \R_DATA_TEMPR28[69] , 
        \R_DATA_TEMPR29[69] , \R_DATA_TEMPR30[69] , 
        \R_DATA_TEMPR31[69] , \R_DATA_TEMPR0[70] , \R_DATA_TEMPR1[70] , 
        \R_DATA_TEMPR2[70] , \R_DATA_TEMPR3[70] , \R_DATA_TEMPR4[70] , 
        \R_DATA_TEMPR5[70] , \R_DATA_TEMPR6[70] , \R_DATA_TEMPR7[70] , 
        \R_DATA_TEMPR8[70] , \R_DATA_TEMPR9[70] , \R_DATA_TEMPR10[70] , 
        \R_DATA_TEMPR11[70] , \R_DATA_TEMPR12[70] , 
        \R_DATA_TEMPR13[70] , \R_DATA_TEMPR14[70] , 
        \R_DATA_TEMPR15[70] , \R_DATA_TEMPR16[70] , 
        \R_DATA_TEMPR17[70] , \R_DATA_TEMPR18[70] , 
        \R_DATA_TEMPR19[70] , \R_DATA_TEMPR20[70] , 
        \R_DATA_TEMPR21[70] , \R_DATA_TEMPR22[70] , 
        \R_DATA_TEMPR23[70] , \R_DATA_TEMPR24[70] , 
        \R_DATA_TEMPR25[70] , \R_DATA_TEMPR26[70] , 
        \R_DATA_TEMPR27[70] , \R_DATA_TEMPR28[70] , 
        \R_DATA_TEMPR29[70] , \R_DATA_TEMPR30[70] , 
        \R_DATA_TEMPR31[70] , \R_DATA_TEMPR0[71] , \R_DATA_TEMPR1[71] , 
        \R_DATA_TEMPR2[71] , \R_DATA_TEMPR3[71] , \R_DATA_TEMPR4[71] , 
        \R_DATA_TEMPR5[71] , \R_DATA_TEMPR6[71] , \R_DATA_TEMPR7[71] , 
        \R_DATA_TEMPR8[71] , \R_DATA_TEMPR9[71] , \R_DATA_TEMPR10[71] , 
        \R_DATA_TEMPR11[71] , \R_DATA_TEMPR12[71] , 
        \R_DATA_TEMPR13[71] , \R_DATA_TEMPR14[71] , 
        \R_DATA_TEMPR15[71] , \R_DATA_TEMPR16[71] , 
        \R_DATA_TEMPR17[71] , \R_DATA_TEMPR18[71] , 
        \R_DATA_TEMPR19[71] , \R_DATA_TEMPR20[71] , 
        \R_DATA_TEMPR21[71] , \R_DATA_TEMPR22[71] , 
        \R_DATA_TEMPR23[71] , \R_DATA_TEMPR24[71] , 
        \R_DATA_TEMPR25[71] , \R_DATA_TEMPR26[71] , 
        \R_DATA_TEMPR27[71] , \R_DATA_TEMPR28[71] , 
        \R_DATA_TEMPR29[71] , \R_DATA_TEMPR30[71] , 
        \R_DATA_TEMPR31[71] , \R_DATA_TEMPR0[72] , \R_DATA_TEMPR1[72] , 
        \R_DATA_TEMPR2[72] , \R_DATA_TEMPR3[72] , \R_DATA_TEMPR4[72] , 
        \R_DATA_TEMPR5[72] , \R_DATA_TEMPR6[72] , \R_DATA_TEMPR7[72] , 
        \R_DATA_TEMPR8[72] , \R_DATA_TEMPR9[72] , \R_DATA_TEMPR10[72] , 
        \R_DATA_TEMPR11[72] , \R_DATA_TEMPR12[72] , 
        \R_DATA_TEMPR13[72] , \R_DATA_TEMPR14[72] , 
        \R_DATA_TEMPR15[72] , \R_DATA_TEMPR16[72] , 
        \R_DATA_TEMPR17[72] , \R_DATA_TEMPR18[72] , 
        \R_DATA_TEMPR19[72] , \R_DATA_TEMPR20[72] , 
        \R_DATA_TEMPR21[72] , \R_DATA_TEMPR22[72] , 
        \R_DATA_TEMPR23[72] , \R_DATA_TEMPR24[72] , 
        \R_DATA_TEMPR25[72] , \R_DATA_TEMPR26[72] , 
        \R_DATA_TEMPR27[72] , \R_DATA_TEMPR28[72] , 
        \R_DATA_TEMPR29[72] , \R_DATA_TEMPR30[72] , 
        \R_DATA_TEMPR31[72] , \R_DATA_TEMPR0[73] , \R_DATA_TEMPR1[73] , 
        \R_DATA_TEMPR2[73] , \R_DATA_TEMPR3[73] , \R_DATA_TEMPR4[73] , 
        \R_DATA_TEMPR5[73] , \R_DATA_TEMPR6[73] , \R_DATA_TEMPR7[73] , 
        \R_DATA_TEMPR8[73] , \R_DATA_TEMPR9[73] , \R_DATA_TEMPR10[73] , 
        \R_DATA_TEMPR11[73] , \R_DATA_TEMPR12[73] , 
        \R_DATA_TEMPR13[73] , \R_DATA_TEMPR14[73] , 
        \R_DATA_TEMPR15[73] , \R_DATA_TEMPR16[73] , 
        \R_DATA_TEMPR17[73] , \R_DATA_TEMPR18[73] , 
        \R_DATA_TEMPR19[73] , \R_DATA_TEMPR20[73] , 
        \R_DATA_TEMPR21[73] , \R_DATA_TEMPR22[73] , 
        \R_DATA_TEMPR23[73] , \R_DATA_TEMPR24[73] , 
        \R_DATA_TEMPR25[73] , \R_DATA_TEMPR26[73] , 
        \R_DATA_TEMPR27[73] , \R_DATA_TEMPR28[73] , 
        \R_DATA_TEMPR29[73] , \R_DATA_TEMPR30[73] , 
        \R_DATA_TEMPR31[73] , \R_DATA_TEMPR0[74] , \R_DATA_TEMPR1[74] , 
        \R_DATA_TEMPR2[74] , \R_DATA_TEMPR3[74] , \R_DATA_TEMPR4[74] , 
        \R_DATA_TEMPR5[74] , \R_DATA_TEMPR6[74] , \R_DATA_TEMPR7[74] , 
        \R_DATA_TEMPR8[74] , \R_DATA_TEMPR9[74] , \R_DATA_TEMPR10[74] , 
        \R_DATA_TEMPR11[74] , \R_DATA_TEMPR12[74] , 
        \R_DATA_TEMPR13[74] , \R_DATA_TEMPR14[74] , 
        \R_DATA_TEMPR15[74] , \R_DATA_TEMPR16[74] , 
        \R_DATA_TEMPR17[74] , \R_DATA_TEMPR18[74] , 
        \R_DATA_TEMPR19[74] , \R_DATA_TEMPR20[74] , 
        \R_DATA_TEMPR21[74] , \R_DATA_TEMPR22[74] , 
        \R_DATA_TEMPR23[74] , \R_DATA_TEMPR24[74] , 
        \R_DATA_TEMPR25[74] , \R_DATA_TEMPR26[74] , 
        \R_DATA_TEMPR27[74] , \R_DATA_TEMPR28[74] , 
        \R_DATA_TEMPR29[74] , \R_DATA_TEMPR30[74] , 
        \R_DATA_TEMPR31[74] , \R_DATA_TEMPR0[75] , \R_DATA_TEMPR1[75] , 
        \R_DATA_TEMPR2[75] , \R_DATA_TEMPR3[75] , \R_DATA_TEMPR4[75] , 
        \R_DATA_TEMPR5[75] , \R_DATA_TEMPR6[75] , \R_DATA_TEMPR7[75] , 
        \R_DATA_TEMPR8[75] , \R_DATA_TEMPR9[75] , \R_DATA_TEMPR10[75] , 
        \R_DATA_TEMPR11[75] , \R_DATA_TEMPR12[75] , 
        \R_DATA_TEMPR13[75] , \R_DATA_TEMPR14[75] , 
        \R_DATA_TEMPR15[75] , \R_DATA_TEMPR16[75] , 
        \R_DATA_TEMPR17[75] , \R_DATA_TEMPR18[75] , 
        \R_DATA_TEMPR19[75] , \R_DATA_TEMPR20[75] , 
        \R_DATA_TEMPR21[75] , \R_DATA_TEMPR22[75] , 
        \R_DATA_TEMPR23[75] , \R_DATA_TEMPR24[75] , 
        \R_DATA_TEMPR25[75] , \R_DATA_TEMPR26[75] , 
        \R_DATA_TEMPR27[75] , \R_DATA_TEMPR28[75] , 
        \R_DATA_TEMPR29[75] , \R_DATA_TEMPR30[75] , 
        \R_DATA_TEMPR31[75] , \R_DATA_TEMPR0[76] , \R_DATA_TEMPR1[76] , 
        \R_DATA_TEMPR2[76] , \R_DATA_TEMPR3[76] , \R_DATA_TEMPR4[76] , 
        \R_DATA_TEMPR5[76] , \R_DATA_TEMPR6[76] , \R_DATA_TEMPR7[76] , 
        \R_DATA_TEMPR8[76] , \R_DATA_TEMPR9[76] , \R_DATA_TEMPR10[76] , 
        \R_DATA_TEMPR11[76] , \R_DATA_TEMPR12[76] , 
        \R_DATA_TEMPR13[76] , \R_DATA_TEMPR14[76] , 
        \R_DATA_TEMPR15[76] , \R_DATA_TEMPR16[76] , 
        \R_DATA_TEMPR17[76] , \R_DATA_TEMPR18[76] , 
        \R_DATA_TEMPR19[76] , \R_DATA_TEMPR20[76] , 
        \R_DATA_TEMPR21[76] , \R_DATA_TEMPR22[76] , 
        \R_DATA_TEMPR23[76] , \R_DATA_TEMPR24[76] , 
        \R_DATA_TEMPR25[76] , \R_DATA_TEMPR26[76] , 
        \R_DATA_TEMPR27[76] , \R_DATA_TEMPR28[76] , 
        \R_DATA_TEMPR29[76] , \R_DATA_TEMPR30[76] , 
        \R_DATA_TEMPR31[76] , \R_DATA_TEMPR0[77] , \R_DATA_TEMPR1[77] , 
        \R_DATA_TEMPR2[77] , \R_DATA_TEMPR3[77] , \R_DATA_TEMPR4[77] , 
        \R_DATA_TEMPR5[77] , \R_DATA_TEMPR6[77] , \R_DATA_TEMPR7[77] , 
        \R_DATA_TEMPR8[77] , \R_DATA_TEMPR9[77] , \R_DATA_TEMPR10[77] , 
        \R_DATA_TEMPR11[77] , \R_DATA_TEMPR12[77] , 
        \R_DATA_TEMPR13[77] , \R_DATA_TEMPR14[77] , 
        \R_DATA_TEMPR15[77] , \R_DATA_TEMPR16[77] , 
        \R_DATA_TEMPR17[77] , \R_DATA_TEMPR18[77] , 
        \R_DATA_TEMPR19[77] , \R_DATA_TEMPR20[77] , 
        \R_DATA_TEMPR21[77] , \R_DATA_TEMPR22[77] , 
        \R_DATA_TEMPR23[77] , \R_DATA_TEMPR24[77] , 
        \R_DATA_TEMPR25[77] , \R_DATA_TEMPR26[77] , 
        \R_DATA_TEMPR27[77] , \R_DATA_TEMPR28[77] , 
        \R_DATA_TEMPR29[77] , \R_DATA_TEMPR30[77] , 
        \R_DATA_TEMPR31[77] , \R_DATA_TEMPR0[78] , \R_DATA_TEMPR1[78] , 
        \R_DATA_TEMPR2[78] , \R_DATA_TEMPR3[78] , \R_DATA_TEMPR4[78] , 
        \R_DATA_TEMPR5[78] , \R_DATA_TEMPR6[78] , \R_DATA_TEMPR7[78] , 
        \R_DATA_TEMPR8[78] , \R_DATA_TEMPR9[78] , \R_DATA_TEMPR10[78] , 
        \R_DATA_TEMPR11[78] , \R_DATA_TEMPR12[78] , 
        \R_DATA_TEMPR13[78] , \R_DATA_TEMPR14[78] , 
        \R_DATA_TEMPR15[78] , \R_DATA_TEMPR16[78] , 
        \R_DATA_TEMPR17[78] , \R_DATA_TEMPR18[78] , 
        \R_DATA_TEMPR19[78] , \R_DATA_TEMPR20[78] , 
        \R_DATA_TEMPR21[78] , \R_DATA_TEMPR22[78] , 
        \R_DATA_TEMPR23[78] , \R_DATA_TEMPR24[78] , 
        \R_DATA_TEMPR25[78] , \R_DATA_TEMPR26[78] , 
        \R_DATA_TEMPR27[78] , \R_DATA_TEMPR28[78] , 
        \R_DATA_TEMPR29[78] , \R_DATA_TEMPR30[78] , 
        \R_DATA_TEMPR31[78] , \R_DATA_TEMPR0[79] , \R_DATA_TEMPR1[79] , 
        \R_DATA_TEMPR2[79] , \R_DATA_TEMPR3[79] , \R_DATA_TEMPR4[79] , 
        \R_DATA_TEMPR5[79] , \R_DATA_TEMPR6[79] , \R_DATA_TEMPR7[79] , 
        \R_DATA_TEMPR8[79] , \R_DATA_TEMPR9[79] , \R_DATA_TEMPR10[79] , 
        \R_DATA_TEMPR11[79] , \R_DATA_TEMPR12[79] , 
        \R_DATA_TEMPR13[79] , \R_DATA_TEMPR14[79] , 
        \R_DATA_TEMPR15[79] , \R_DATA_TEMPR16[79] , 
        \R_DATA_TEMPR17[79] , \R_DATA_TEMPR18[79] , 
        \R_DATA_TEMPR19[79] , \R_DATA_TEMPR20[79] , 
        \R_DATA_TEMPR21[79] , \R_DATA_TEMPR22[79] , 
        \R_DATA_TEMPR23[79] , \R_DATA_TEMPR24[79] , 
        \R_DATA_TEMPR25[79] , \R_DATA_TEMPR26[79] , 
        \R_DATA_TEMPR27[79] , \R_DATA_TEMPR28[79] , 
        \R_DATA_TEMPR29[79] , \R_DATA_TEMPR30[79] , 
        \R_DATA_TEMPR31[79] , \BLKX0[0] , \BLKY0[0] , \BLKX1[0] , 
        \BLKY1[0] , \BLKX2[0] , \BLKX2[1] , \BLKX2[2] , \BLKX2[3] , 
        \BLKX2[4] , \BLKX2[5] , \BLKX2[6] , \BLKX2[7] , \BLKY2[0] , 
        \BLKY2[1] , \BLKY2[2] , \BLKY2[3] , \BLKY2[4] , \BLKY2[5] , 
        \BLKY2[6] , \BLKY2[7] , \ACCESS_BUSY[0][0] , 
        \ACCESS_BUSY[0][1] , \ACCESS_BUSY[1][0] , \ACCESS_BUSY[1][1] , 
        \ACCESS_BUSY[2][0] , \ACCESS_BUSY[2][1] , \ACCESS_BUSY[3][0] , 
        \ACCESS_BUSY[3][1] , \ACCESS_BUSY[4][0] , \ACCESS_BUSY[4][1] , 
        \ACCESS_BUSY[5][0] , \ACCESS_BUSY[5][1] , \ACCESS_BUSY[6][0] , 
        \ACCESS_BUSY[6][1] , \ACCESS_BUSY[7][0] , \ACCESS_BUSY[7][1] , 
        \ACCESS_BUSY[8][0] , \ACCESS_BUSY[8][1] , \ACCESS_BUSY[9][0] , 
        \ACCESS_BUSY[9][1] , \ACCESS_BUSY[10][0] , 
        \ACCESS_BUSY[10][1] , \ACCESS_BUSY[11][0] , 
        \ACCESS_BUSY[11][1] , \ACCESS_BUSY[12][0] , 
        \ACCESS_BUSY[12][1] , \ACCESS_BUSY[13][0] , 
        \ACCESS_BUSY[13][1] , \ACCESS_BUSY[14][0] , 
        \ACCESS_BUSY[14][1] , \ACCESS_BUSY[15][0] , 
        \ACCESS_BUSY[15][1] , \ACCESS_BUSY[16][0] , 
        \ACCESS_BUSY[16][1] , \ACCESS_BUSY[17][0] , 
        \ACCESS_BUSY[17][1] , \ACCESS_BUSY[18][0] , 
        \ACCESS_BUSY[18][1] , \ACCESS_BUSY[19][0] , 
        \ACCESS_BUSY[19][1] , \ACCESS_BUSY[20][0] , 
        \ACCESS_BUSY[20][1] , \ACCESS_BUSY[21][0] , 
        \ACCESS_BUSY[21][1] , \ACCESS_BUSY[22][0] , 
        \ACCESS_BUSY[22][1] , \ACCESS_BUSY[23][0] , 
        \ACCESS_BUSY[23][1] , \ACCESS_BUSY[24][0] , 
        \ACCESS_BUSY[24][1] , \ACCESS_BUSY[25][0] , 
        \ACCESS_BUSY[25][1] , \ACCESS_BUSY[26][0] , 
        \ACCESS_BUSY[26][1] , \ACCESS_BUSY[27][0] , 
        \ACCESS_BUSY[27][1] , \ACCESS_BUSY[28][0] , 
        \ACCESS_BUSY[28][1] , \ACCESS_BUSY[29][0] , 
        \ACCESS_BUSY[29][1] , \ACCESS_BUSY[30][0] , 
        \ACCESS_BUSY[30][1] , \ACCESS_BUSY[31][0] , 
        \ACCESS_BUSY[31][1] , CFG2_3_Y, CFG2_6_Y, CFG2_1_Y, CFG2_5_Y, 
        OR4_392_Y, OR4_358_Y, OR4_499_Y, OR4_551_Y, OR4_474_Y, 
        OR4_231_Y, OR4_478_Y, OR4_215_Y, OR4_490_Y, OR2_46_Y, OR4_87_Y, 
        OR4_433_Y, OR4_624_Y, OR4_692_Y, OR4_151_Y, OR4_554_Y, 
        OR4_98_Y, OR4_450_Y, OR4_331_Y, OR2_71_Y, OR4_37_Y, OR4_214_Y, 
        OR4_529_Y, OR4_264_Y, OR4_703_Y, OR4_549_Y, OR4_711_Y, 
        OR4_311_Y, OR4_306_Y, OR2_25_Y, OR4_700_Y, OR4_664_Y, 
        OR4_674_Y, OR4_447_Y, OR4_229_Y, OR4_342_Y, OR4_337_Y, 
        OR4_455_Y, OR4_150_Y, OR2_3_Y, OR4_256_Y, OR4_403_Y, OR4_10_Y, 
        OR4_454_Y, OR4_199_Y, OR4_35_Y, OR4_207_Y, OR4_523_Y, 
        OR4_518_Y, OR2_5_Y, OR4_611_Y, OR4_419_Y, OR4_391_Y, OR4_366_Y, 
        OR4_116_Y, OR4_709_Y, OR4_693_Y, OR4_409_Y, OR4_285_Y, OR2_6_Y, 
        OR4_88_Y, OR4_628_Y, OR4_603_Y, OR4_577_Y, OR4_325_Y, 
        OR4_201_Y, OR4_185_Y, OR4_620_Y, OR4_496_Y, OR2_70_Y, 
        OR4_131_Y, OR4_300_Y, OR4_632_Y, OR4_349_Y, OR4_72_Y, 
        OR4_651_Y, OR4_79_Y, OR4_414_Y, OR4_406_Y, OR2_11_Y, OR4_178_Y, 
        OR4_373_Y, OR4_314_Y, OR4_371_Y, OR4_224_Y, OR4_453_Y, 
        OR4_642_Y, OR4_254_Y, OR4_293_Y, OR2_21_Y, OR4_189_Y, 
        OR4_652_Y, OR4_283_Y, OR4_598_Y, OR4_59_Y, OR4_226_Y, 
        OR4_295_Y, OR4_93_Y, OR4_112_Y, OR2_60_Y, OR4_712_Y, OR4_521_Y, 
        OR4_493_Y, OR4_470_Y, OR4_238_Y, OR4_75_Y, OR4_64_Y, OR4_514_Y, 
        OR4_389_Y, OR2_75_Y, OR4_125_Y, OR4_38_Y, OR4_425_Y, OR4_531_Y, 
        OR4_638_Y, OR4_488_Y, OR4_365_Y, OR4_396_Y, OR4_377_Y, 
        OR2_37_Y, OR4_338_Y, OR4_258_Y, OR4_641_Y, OR4_13_Y, OR4_111_Y, 
        OR4_694_Y, OR4_574_Y, OR4_609_Y, OR4_587_Y, OR2_16_Y, 
        OR4_362_Y, OR4_441_Y, OR4_275_Y, OR4_542_Y, OR4_100_Y, 
        OR4_149_Y, OR4_387_Y, OR4_143_Y, OR4_479_Y, OR2_42_Y, 
        OR4_249_Y, OR4_133_Y, OR4_532_Y, OR4_634_Y, OR4_12_Y, 
        OR4_588_Y, OR4_465_Y, OR4_500_Y, OR4_483_Y, OR2_27_Y, 
        OR4_280_Y, OR4_673_Y, OR4_68_Y, OR4_101_Y, OR4_629_Y, 
        OR4_407_Y, OR4_446_Y, OR4_579_Y, OR4_104_Y, OR2_9_Y, OR4_171_Y, 
        OR4_9_Y, OR4_681_Y, OR4_561_Y, OR4_458_Y, OR4_704_Y, OR4_288_Y, 
        OR4_585_Y, OR4_319_Y, OR2_79_Y, OR4_107_Y, OR4_688_Y, 
        OR4_457_Y, OR4_601_Y, OR4_321_Y, OR4_575_Y, OR4_516_Y, 
        OR4_228_Y, OR4_105_Y, OR2_13_Y, OR4_170_Y, OR4_126_Y, 
        OR4_142_Y, OR4_648_Y, OR4_415_Y, OR4_540_Y, OR4_538_Y, 
        OR4_653_Y, OR4_345_Y, OR2_39_Y, OR4_462_Y, OR4_437_Y, 
        OR4_339_Y, OR4_18_Y, OR4_596_Y, OR4_297_Y, OR4_445_Y, OR4_80_Y, 
        OR4_128_Y, OR2_35_Y, OR4_378_Y, OR4_341_Y, OR4_352_Y, 
        OR4_120_Y, OR4_623_Y, OR4_23_Y, OR4_22_Y, OR4_135_Y, OR4_559_Y, 
        OR2_22_Y, OR4_154_Y, OR4_501_Y, OR4_682_Y, OR4_29_Y, OR4_223_Y, 
        OR4_614_Y, OR4_167_Y, OR4_512_Y, OR4_397_Y, OR2_47_Y, 
        OR4_277_Y, OR4_250_Y, OR4_261_Y, OR4_25_Y, OR4_517_Y, 
        OR4_643_Y, OR4_640_Y, OR4_33_Y, OR4_442_Y, OR2_31_Y, OR4_81_Y, 
        OR4_263_Y, OR4_578_Y, OR4_299_Y, OR4_30_Y, OR4_600_Y, OR4_36_Y, 
        OR4_364_Y, OR4_355_Y, OR2_50_Y, OR4_571_Y, OR4_205_Y, 
        OR4_472_Y, OR4_274_Y, OR4_123_Y, OR4_552_Y, OR4_582_Y, 
        OR4_237_Y, OR4_637_Y, OR2_44_Y, OR4_658_Y, OR4_469_Y, 
        OR4_435_Y, OR4_420_Y, OR4_184_Y, OR4_31_Y, OR4_21_Y, OR4_460_Y, 
        OR4_333_Y, OR2_34_Y, OR4_422_Y, OR4_661_Y, OR4_459_Y, 
        OR4_353_Y, OR4_696_Y, OR4_96_Y, OR4_533_Y, OR4_443_Y, 
        OR4_211_Y, OR2_49_Y, OR4_191_Y, OR4_83_Y, OR4_482_Y, OR4_580_Y, 
        OR4_683_Y, OR4_537_Y, OR4_413_Y, OR4_444_Y, OR4_424_Y, 
        OR2_61_Y, OR4_330_Y, OR4_6_Y, OR4_129_Y, OR4_173_Y, OR4_684_Y, 
        OR4_471_Y, OR4_509_Y, OR4_645_Y, OR4_182_Y, OR2_67_Y, 
        OR4_240_Y, OR4_66_Y, OR4_24_Y, OR4_621_Y, OR4_524_Y, OR4_40_Y, 
        OR4_347_Y, OR4_649_Y, OR4_386_Y, OR2_55_Y, CFG2_4_Y, CFG2_2_Y, 
        CFG2_7_Y, CFG2_0_Y, OR4_589_Y, OR4_677_Y, OR4_480_Y, OR4_384_Y, 
        OR4_665_Y, OR4_11_Y, OR4_63_Y, OR4_16_Y, OR4_427_Y, OR2_68_Y, 
        OR4_526_Y, OR4_502_Y, OR4_398_Y, OR4_69_Y, OR4_656_Y, 
        OR4_356_Y, OR4_508_Y, OR4_144_Y, OR4_209_Y, OR2_4_Y, OR4_117_Y, 
        OR4_473_Y, OR4_657_Y, OR4_717_Y, OR4_195_Y, OR4_584_Y, 
        OR4_137_Y, OR4_489_Y, OR4_370_Y, OR2_23_Y, OR4_230_Y, 
        OR4_193_Y, OR4_210_Y, OR4_697_Y, OR4_464_Y, OR4_590_Y, 
        OR4_586_Y, OR4_710_Y, OR4_394_Y, OR2_63_Y, OR4_636_Y, 
        OR4_265_Y, OR4_535_Y, OR4_320_Y, OR4_204_Y, OR4_612_Y, 
        OR4_646_Y, OR4_284_Y, OR4_695_Y, OR2_18_Y, OR4_630_Y, 
        OR4_374_Y, OR4_4_Y, OR4_315_Y, OR4_511_Y, OR4_666_Y, OR4_20_Y, 
        OR4_550_Y, OR4_569_Y, OR2_51_Y, OR4_309_Y, OR4_705_Y, OR4_97_Y, 
        OR4_141_Y, OR4_659_Y, OR4_438_Y, OR4_487_Y, OR4_613_Y, 
        OR4_146_Y, OR2_43_Y, OR4_90_Y, OR4_242_Y, OR4_417_Y, OR4_560_Y, 
        OR4_239_Y, OR4_639_Y, OR4_399_Y, OR4_157_Y, OR4_375_Y, 
        OR2_10_Y, OR4_218_Y, OR4_42_Y, OR4_714_Y, OR4_595_Y, OR4_492_Y, 
        OR4_7_Y, OR4_318_Y, OR4_617_Y, OR4_357_Y, OR2_33_Y, OR4_316_Y, 
        OR4_670_Y, OR4_119_Y, OR4_208_Y, OR4_379_Y, OR4_53_Y, 
        OR4_328_Y, OR4_678_Y, OR4_563_Y, OR2_58_Y, OR4_530_Y, 
        OR4_153_Y, OR4_329_Y, OR4_400_Y, OR4_591_Y, OR4_273_Y, 
        OR4_545_Y, OR4_162_Y, OR4_46_Y, OR2_38_Y, OR4_495_Y, OR4_476_Y, 
        OR4_372_Y, OR4_45_Y, OR4_626_Y, OR4_322_Y, OR4_486_Y, 
        OR4_108_Y, OR4_165_Y, OR2_64_Y, OR4_421_Y, OR4_43_Y, OR4_241_Y, 
        OR4_294_Y, OR4_484_Y, OR4_158_Y, OR4_429_Y, OR4_55_Y, 
        OR4_668_Y, OR2_45_Y, OR4_599_Y, OR4_680_Y, OR4_452_Y, 
        OR4_592_Y, OR4_573_Y, OR4_568_Y, OR4_525_Y, OR4_702_Y, 
        OR4_99_Y, OR2_69_Y, OR4_605_Y, OR4_234_Y, OR4_505_Y, OR4_298_Y, 
        OR4_161_Y, OR4_583_Y, OR4_615_Y, OR4_269_Y, OR4_667_Y, 
        OR2_73_Y, OR4_534_Y, OR4_698_Y, OR4_301_Y, OR4_26_Y, OR4_475_Y, 
        OR4_317_Y, OR4_485_Y, OR4_82_Y, OR4_74_Y, OR2_40_Y, OR4_383_Y, 
        OR4_206_Y, OR4_164_Y, OR4_139_Y, OR4_622_Y, OR4_477_Y, 
        OR4_466_Y, OR4_197_Y, OR4_57_Y, OR2_24_Y, OR4_504_Y, OR4_176_Y, 
        OR4_302_Y, OR4_332_Y, OR4_121_Y, OR4_644_Y, OR4_676_Y, 
        OR4_73_Y, OR4_340_Y, OR2_74_Y, OR4_686_Y, OR4_428_Y, OR4_60_Y, 
        OR4_380_Y, OR4_572_Y, OR4_718_Y, OR4_71_Y, OR4_610_Y, 
        OR4_631_Y, OR2_28_Y, OR4_713_Y, OR4_381_Y, OR4_510_Y, 
        OR4_548_Y, OR4_334_Y, OR4_114_Y, OR4_160_Y, OR4_287_Y, 
        OR4_553_Y, OR2_59_Y, OR4_393_Y, OR4_252_Y, OR4_202_Y, OR4_58_Y, 
        OR4_685_Y, OR4_221_Y, OR4_519_Y, OR4_85_Y, OR4_555_Y, OR2_65_Y, 
        OR4_607_Y, OR4_440_Y, OR4_395_Y, OR4_278_Y, OR4_177_Y, 
        OR4_410_Y, OR4_719_Y, OR4_296_Y, OR4_41_Y, OR2_48_Y, OR4_633_Y, 
        OR4_536_Y, OR4_217_Y, OR4_303_Y, OR4_405_Y, OR4_268_Y, 
        OR4_132_Y, OR4_172_Y, OR4_148_Y, OR2_52_Y, OR4_608_Y, 
        OR4_279_Y, OR4_401_Y, OR4_431_Y, OR4_245_Y, OR4_17_Y, OR4_52_Y, 
        OR4_192_Y, OR4_436_Y, OR2_66_Y, OR4_497_Y, OR4_336_Y, 
        OR4_290_Y, OR4_163_Y, OR4_61_Y, OR4_304_Y, OR4_619_Y, 
        OR4_203_Y, OR4_655_Y, OR2_54_Y, OR4_690_Y, OR4_672_Y, 
        OR4_567_Y, OR4_255_Y, OR4_91_Y, OR4_527_Y, OR4_675_Y, 
        OR4_310_Y, OR4_360_Y, OR2_14_Y, OR4_183_Y, OR4_156_Y, OR4_49_Y, 
        OR4_448_Y, OR4_305_Y, OR4_8_Y, OR4_159_Y, OR4_522_Y, OR4_570_Y, 
        OR2_77_Y, OR4_168_Y, OR4_515_Y, OR4_27_Y, OR4_118_Y, OR4_92_Y, 
        OR4_327_Y, OR4_179_Y, OR4_174_Y, OR4_140_Y, OR2_19_Y, 
        OR4_369_Y, OR4_715_Y, OR4_186_Y, OR4_257_Y, OR4_426_Y, 
        OR4_95_Y, OR4_385_Y, OR4_5_Y, OR4_616_Y, OR2_78_Y, OR4_62_Y, 
        OR4_44_Y, OR4_671_Y, OR4_344_Y, OR4_216_Y, OR4_625_Y, OR4_51_Y, 
        OR4_411_Y, OR4_461_Y, OR2_2_Y, OR4_67_Y, OR4_418_Y, OR4_701_Y, 
        OR4_494_Y, OR4_354_Y, OR4_50_Y, OR4_77_Y, OR4_449_Y, OR4_130_Y, 
        OR2_30_Y, OR4_282_Y, OR4_627_Y, OR4_194_Y, OR4_707_Y, 
        OR4_565_Y, OR4_271_Y, OR4_291_Y, OR4_663_Y, OR4_343_Y, OR2_8_Y, 
        OR4_669_Y, OR4_635_Y, OR4_647_Y, OR4_416_Y, OR4_200_Y, 
        OR4_308_Y, OR4_307_Y, OR4_423_Y, OR4_110_Y, OR2_56_Y, 
        OR4_181_Y, OR4_520_Y, OR4_70_Y, OR4_597_Y, OR4_456_Y, 
        OR4_155_Y, OR4_196_Y, OR4_557_Y, OR4_251_Y, OR2_17_Y, 
        OR4_593_Y, OR4_34_Y, OR4_359_Y, OR4_76_Y, OR4_539_Y, OR4_382_Y, 
        OR4_543_Y, OR4_145_Y, OR4_138_Y, OR2_12_Y, OR4_556_Y, 
        OR4_136_Y, OR4_246_Y, OR4_312_Y, OR4_78_Y, OR4_225_Y, OR4_86_Y, 
        OR4_463_Y, OR4_56_Y, OR2_62_Y, OR4_434_Y, OR4_266_Y, OR4_236_Y, 
        OR4_219_Y, OR4_679_Y, OR4_541_Y, OR4_528_Y, OR4_260_Y, 
        OR4_113_Y, OR2_76_Y, OR4_660_Y, OR4_402_Y, OR4_39_Y, OR4_348_Y, 
        OR4_544_Y, OR4_699_Y, OR4_48_Y, OR4_581_Y, OR4_602_Y, OR2_0_Y, 
        OR4_558_Y, OR4_233_Y, OR4_350_Y, OR4_388_Y, OR4_188_Y, 
        OR4_687_Y, OR4_1_Y, OR4_124_Y, OR4_390_Y, OR2_20_Y, OR4_439_Y, 
        OR4_286_Y, OR4_253_Y, OR4_103_Y, OR4_15_Y, OR4_267_Y, 
        OR4_566_Y, OR4_134_Y, OR4_606_Y, OR2_7_Y, OR4_689_Y, OR4_594_Y, 
        OR4_272_Y, OR4_361_Y, OR4_467_Y, OR4_313_Y, OR4_212_Y, 
        OR4_244_Y, OR4_222_Y, OR2_29_Y, OR4_19_Y, OR4_716_Y, OR4_618_Y, 
        OR4_292_Y, OR4_147_Y, OR4_576_Y, OR4_0_Y, OR4_363_Y, OR4_408_Y, 
        OR2_41_Y, OR4_115_Y, OR4_468_Y, OR4_28_Y, OR4_546_Y, OR4_404_Y, 
        OR4_94_Y, OR4_127_Y, OR4_503_Y, OR4_198_Y, OR2_53_Y, OR4_2_Y, 
        OR4_691_Y, OR4_706_Y, OR4_481_Y, OR4_262_Y, OR4_368_Y, 
        OR4_367_Y, OR4_491_Y, OR4_187_Y, OR2_32_Y, OR4_562_Y, OR4_3_Y, 
        OR4_323_Y, OR4_54_Y, OR4_506_Y, OR4_351_Y, OR4_513_Y, 
        OR4_109_Y, OR4_102_Y, OR2_72_Y, OR4_122_Y, OR4_604_Y, 
        OR4_243_Y, OR4_547_Y, OR4_14_Y, OR4_166_Y, OR4_259_Y, OR4_47_Y, 
        OR4_65_Y, OR2_36_Y, OR4_335_Y, OR4_84_Y, OR4_430_Y, OR4_32_Y, 
        OR4_232_Y, OR4_376_Y, OR4_451_Y, OR4_270_Y, OR4_281_Y, 
        OR2_15_Y, OR4_412_Y, OR4_235_Y, OR4_213_Y, OR4_180_Y, 
        OR4_654_Y, OR4_507_Y, OR4_498_Y, OR4_227_Y, OR4_89_Y, OR2_57_Y, 
        OR4_247_Y, OR4_708_Y, OR4_324_Y, OR4_650_Y, OR4_106_Y, 
        OR4_276_Y, OR4_346_Y, OR4_152_Y, OR4_175_Y, OR2_26_Y, 
        OR4_662_Y, OR4_564_Y, OR4_248_Y, OR4_326_Y, OR4_432_Y, 
        OR4_289_Y, OR4_169_Y, OR4_220_Y, OR4_190_Y, OR2_1_Y, VCC, GND, 
        ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    OR4 OR4_700 (.A(OR4_229_Y), .B(OR4_342_Y), .C(OR4_337_Y), .D(
        OR4_455_Y), .Y(OR4_700_Y));
    OR4 OR4_399 (.A(\R_DATA_TEMPR8[9] ), .B(\R_DATA_TEMPR9[9] ), .C(
        \R_DATA_TEMPR10[9] ), .D(\R_DATA_TEMPR11[9] ), .Y(OR4_399_Y));
    OR4 OR4_420 (.A(\R_DATA_TEMPR28[63] ), .B(\R_DATA_TEMPR29[63] ), 
        .C(\R_DATA_TEMPR30[63] ), .D(\R_DATA_TEMPR31[63] ), .Y(
        OR4_420_Y));
    OR4 OR4_402 (.A(OR4_602_Y), .B(OR2_0_Y), .C(\R_DATA_TEMPR22[74] ), 
        .D(\R_DATA_TEMPR23[74] ), .Y(OR4_402_Y));
    OR4 OR4_384 (.A(\R_DATA_TEMPR28[1] ), .B(\R_DATA_TEMPR29[1] ), .C(
        \R_DATA_TEMPR30[1] ), .D(\R_DATA_TEMPR31[1] ), .Y(OR4_384_Y));
    OR4 OR4_373 (.A(OR4_293_Y), .B(OR2_21_Y), .C(\R_DATA_TEMPR22[3] ), 
        .D(\R_DATA_TEMPR23[3] ), .Y(OR4_373_Y));
    OR4 \OR4_R_DATA[59]  (.A(OR4_497_Y), .B(OR4_336_Y), .C(OR4_290_Y), 
        .D(OR4_163_Y), .Y(R_DATA[59]));
    OR4 OR4_253 (.A(\R_DATA_TEMPR24[69] ), .B(\R_DATA_TEMPR25[69] ), 
        .C(\R_DATA_TEMPR26[69] ), .D(\R_DATA_TEMPR27[69] ), .Y(
        OR4_253_Y));
    OR4 OR4_409 (.A(\R_DATA_TEMPR12[33] ), .B(\R_DATA_TEMPR13[33] ), 
        .C(\R_DATA_TEMPR14[33] ), .D(\R_DATA_TEMPR15[33] ), .Y(
        OR4_409_Y));
    OR4 OR4_472 (.A(\R_DATA_TEMPR24[25] ), .B(\R_DATA_TEMPR25[25] ), 
        .C(\R_DATA_TEMPR26[25] ), .D(\R_DATA_TEMPR27[25] ), .Y(
        OR4_472_Y));
    OR4 OR4_181 (.A(OR4_456_Y), .B(OR4_155_Y), .C(OR4_196_Y), .D(
        OR4_557_Y), .Y(OR4_181_Y));
    OR4 OR4_106 (.A(\R_DATA_TEMPR0[54] ), .B(\R_DATA_TEMPR1[54] ), .C(
        \R_DATA_TEMPR2[54] ), .D(\R_DATA_TEMPR3[54] ), .Y(OR4_106_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[2]  (.A(CFG2_7_Y), .B(
        W_ADDR[13]), .C(W_EN), .Y(\BLKX2[2] ));
    OR4 OR4_83 (.A(OR4_424_Y), .B(OR2_61_Y), .C(\R_DATA_TEMPR22[68] ), 
        .D(\R_DATA_TEMPR23[68] ), .Y(OR4_83_Y));
    OR4 OR4_479 (.A(\R_DATA_TEMPR16[8] ), .B(\R_DATA_TEMPR17[8] ), .C(
        \R_DATA_TEMPR18[8] ), .D(\R_DATA_TEMPR19[8] ), .Y(OR4_479_Y));
    OR4 OR4_138 (.A(\R_DATA_TEMPR16[10] ), .B(\R_DATA_TEMPR17[10] ), 
        .C(\R_DATA_TEMPR18[10] ), .D(\R_DATA_TEMPR19[10] ), .Y(
        OR4_138_Y));
    OR4 OR4_176 (.A(OR4_340_Y), .B(OR2_74_Y), .C(\R_DATA_TEMPR22[36] ), 
        .D(\R_DATA_TEMPR23[36] ), .Y(OR4_176_Y));
    OR4 OR4_610 (.A(\R_DATA_TEMPR12[14] ), .B(\R_DATA_TEMPR13[14] ), 
        .C(\R_DATA_TEMPR14[14] ), .D(\R_DATA_TEMPR15[14] ), .Y(
        OR4_610_Y));
    OR2 OR2_43 (.A(\R_DATA_TEMPR20[76] ), .B(\R_DATA_TEMPR21[76] ), .Y(
        OR2_43_Y));
    OR4 OR4_481 (.A(\R_DATA_TEMPR28[11] ), .B(\R_DATA_TEMPR29[11] ), 
        .C(\R_DATA_TEMPR30[11] ), .D(\R_DATA_TEMPR31[11] ), .Y(
        OR4_481_Y));
    OR4 OR4_488 (.A(\R_DATA_TEMPR4[38] ), .B(\R_DATA_TEMPR5[38] ), .C(
        \R_DATA_TEMPR6[38] ), .D(\R_DATA_TEMPR7[38] ), .Y(OR4_488_Y));
    OR4 OR4_308 (.A(\R_DATA_TEMPR4[21] ), .B(\R_DATA_TEMPR5[21] ), .C(
        \R_DATA_TEMPR6[21] ), .D(\R_DATA_TEMPR7[21] ), .Y(OR4_308_Y));
    OR4 OR4_317 (.A(\R_DATA_TEMPR4[20] ), .B(\R_DATA_TEMPR5[20] ), .C(
        \R_DATA_TEMPR6[20] ), .D(\R_DATA_TEMPR7[20] ), .Y(OR4_317_Y));
    OR4 OR4_110 (.A(\R_DATA_TEMPR16[21] ), .B(\R_DATA_TEMPR17[21] ), 
        .C(\R_DATA_TEMPR18[21] ), .D(\R_DATA_TEMPR19[21] ), .Y(
        OR4_110_Y));
    OR4 OR4_658 (.A(OR4_184_Y), .B(OR4_31_Y), .C(OR4_21_Y), .D(
        OR4_460_Y), .Y(OR4_658_Y));
    OR4 OR4_378 (.A(OR4_623_Y), .B(OR4_23_Y), .C(OR4_22_Y), .D(
        OR4_135_Y), .Y(OR4_378_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%2%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C1 (
        .A_DOUT({\R_DATA_TEMPR2[79] , \R_DATA_TEMPR2[78] , 
        \R_DATA_TEMPR2[77] , \R_DATA_TEMPR2[76] , \R_DATA_TEMPR2[75] , 
        \R_DATA_TEMPR2[74] , \R_DATA_TEMPR2[73] , \R_DATA_TEMPR2[72] , 
        \R_DATA_TEMPR2[71] , \R_DATA_TEMPR2[70] , \R_DATA_TEMPR2[69] , 
        \R_DATA_TEMPR2[68] , \R_DATA_TEMPR2[67] , \R_DATA_TEMPR2[66] , 
        \R_DATA_TEMPR2[65] , \R_DATA_TEMPR2[64] , \R_DATA_TEMPR2[63] , 
        \R_DATA_TEMPR2[62] , \R_DATA_TEMPR2[61] , \R_DATA_TEMPR2[60] })
        , .B_DOUT({\R_DATA_TEMPR2[59] , \R_DATA_TEMPR2[58] , 
        \R_DATA_TEMPR2[57] , \R_DATA_TEMPR2[56] , \R_DATA_TEMPR2[55] , 
        \R_DATA_TEMPR2[54] , \R_DATA_TEMPR2[53] , \R_DATA_TEMPR2[52] , 
        \R_DATA_TEMPR2[51] , \R_DATA_TEMPR2[50] , \R_DATA_TEMPR2[49] , 
        \R_DATA_TEMPR2[48] , \R_DATA_TEMPR2[47] , \R_DATA_TEMPR2[46] , 
        \R_DATA_TEMPR2[45] , \R_DATA_TEMPR2[44] , \R_DATA_TEMPR2[43] , 
        \R_DATA_TEMPR2[42] , \R_DATA_TEMPR2[41] , \R_DATA_TEMPR2[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[2][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[0] , 
        R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[0] , W_ADDR[10], \BLKX0[0] }), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_2 (.A(OR4_262_Y), .B(OR4_368_Y), .C(OR4_367_Y), .D(
        OR4_491_Y), .Y(OR4_2_Y));
    OR4 OR4_718 (.A(\R_DATA_TEMPR4[14] ), .B(\R_DATA_TEMPR5[14] ), .C(
        \R_DATA_TEMPR6[14] ), .D(\R_DATA_TEMPR7[14] ), .Y(OR4_718_Y));
    OR2 OR2_75 (.A(\R_DATA_TEMPR20[53] ), .B(\R_DATA_TEMPR21[53] ), .Y(
        OR2_75_Y));
    OR4 OR4_329 (.A(\R_DATA_TEMPR24[47] ), .B(\R_DATA_TEMPR25[47] ), 
        .C(\R_DATA_TEMPR26[47] ), .D(\R_DATA_TEMPR27[47] ), .Y(
        OR4_329_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%22%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C1 (
        .A_DOUT({\R_DATA_TEMPR22[79] , \R_DATA_TEMPR22[78] , 
        \R_DATA_TEMPR22[77] , \R_DATA_TEMPR22[76] , 
        \R_DATA_TEMPR22[75] , \R_DATA_TEMPR22[74] , 
        \R_DATA_TEMPR22[73] , \R_DATA_TEMPR22[72] , 
        \R_DATA_TEMPR22[71] , \R_DATA_TEMPR22[70] , 
        \R_DATA_TEMPR22[69] , \R_DATA_TEMPR22[68] , 
        \R_DATA_TEMPR22[67] , \R_DATA_TEMPR22[66] , 
        \R_DATA_TEMPR22[65] , \R_DATA_TEMPR22[64] , 
        \R_DATA_TEMPR22[63] , \R_DATA_TEMPR22[62] , 
        \R_DATA_TEMPR22[61] , \R_DATA_TEMPR22[60] }), .B_DOUT({
        \R_DATA_TEMPR22[59] , \R_DATA_TEMPR22[58] , 
        \R_DATA_TEMPR22[57] , \R_DATA_TEMPR22[56] , 
        \R_DATA_TEMPR22[55] , \R_DATA_TEMPR22[54] , 
        \R_DATA_TEMPR22[53] , \R_DATA_TEMPR22[52] , 
        \R_DATA_TEMPR22[51] , \R_DATA_TEMPR22[50] , 
        \R_DATA_TEMPR22[49] , \R_DATA_TEMPR22[48] , 
        \R_DATA_TEMPR22[47] , \R_DATA_TEMPR22[46] , 
        \R_DATA_TEMPR22[45] , \R_DATA_TEMPR22[44] , 
        \R_DATA_TEMPR22[43] , \R_DATA_TEMPR22[42] , 
        \R_DATA_TEMPR22[41] , \R_DATA_TEMPR22[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[22][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[29]  (.A(OR4_171_Y), .B(OR4_9_Y), .C(OR4_681_Y), 
        .D(OR4_561_Y), .Y(R_DATA[29]));
    OR2 OR2_63 (.A(\R_DATA_TEMPR20[61] ), .B(\R_DATA_TEMPR21[61] ), .Y(
        OR2_63_Y));
    OR4 OR4_667 (.A(\R_DATA_TEMPR16[75] ), .B(\R_DATA_TEMPR17[75] ), 
        .C(\R_DATA_TEMPR18[75] ), .D(\R_DATA_TEMPR19[75] ), .Y(
        OR4_667_Y));
    OR4 OR4_652 (.A(OR4_112_Y), .B(OR2_60_Y), .C(\R_DATA_TEMPR22[64] ), 
        .D(\R_DATA_TEMPR23[64] ), .Y(OR4_652_Y));
    OR4 OR4_593 (.A(OR4_539_Y), .B(OR4_382_Y), .C(OR4_543_Y), .D(
        OR4_145_Y), .Y(OR4_593_Y));
    OR4 OR4_48 (.A(\R_DATA_TEMPR8[74] ), .B(\R_DATA_TEMPR9[74] ), .C(
        \R_DATA_TEMPR10[74] ), .D(\R_DATA_TEMPR11[74] ), .Y(OR4_48_Y));
    OR4 OR4_589 (.A(OR4_665_Y), .B(OR4_11_Y), .C(OR4_63_Y), .D(
        OR4_16_Y), .Y(OR4_589_Y));
    OR4 OR4_109 (.A(\R_DATA_TEMPR12[70] ), .B(\R_DATA_TEMPR13[70] ), 
        .C(\R_DATA_TEMPR14[70] ), .D(\R_DATA_TEMPR15[70] ), .Y(
        OR4_109_Y));
    OR2 OR2_33 (.A(\R_DATA_TEMPR20[79] ), .B(\R_DATA_TEMPR21[79] ), .Y(
        OR2_33_Y));
    OR2 OR2_15 (.A(\R_DATA_TEMPR20[44] ), .B(\R_DATA_TEMPR21[44] ), .Y(
        OR2_15_Y));
    OR4 OR4_241 (.A(\R_DATA_TEMPR24[57] ), .B(\R_DATA_TEMPR25[57] ), 
        .C(\R_DATA_TEMPR26[57] ), .D(\R_DATA_TEMPR27[57] ), .Y(
        OR4_241_Y));
    OR4 OR4_580 (.A(\R_DATA_TEMPR28[68] ), .B(\R_DATA_TEMPR29[68] ), 
        .C(\R_DATA_TEMPR30[68] ), .D(\R_DATA_TEMPR31[68] ), .Y(
        OR4_580_Y));
    OR4 OR4_81 (.A(OR4_30_Y), .B(OR4_600_Y), .C(OR4_36_Y), .D(
        OR4_364_Y), .Y(OR4_81_Y));
    OR4 OR4_118 (.A(\R_DATA_TEMPR28[6] ), .B(\R_DATA_TEMPR29[6] ), .C(
        \R_DATA_TEMPR30[6] ), .D(\R_DATA_TEMPR31[6] ), .Y(OR4_118_Y));
    OR4 \OR4_R_DATA[7]  (.A(OR4_422_Y), .B(OR4_661_Y), .C(OR4_459_Y), 
        .D(OR4_353_Y), .Y(R_DATA[7]));
    OR4 OR4_179 (.A(\R_DATA_TEMPR8[6] ), .B(\R_DATA_TEMPR9[6] ), .C(
        \R_DATA_TEMPR10[6] ), .D(\R_DATA_TEMPR11[6] ), .Y(OR4_179_Y));
    OR2 OR2_41 (.A(\R_DATA_TEMPR20[62] ), .B(\R_DATA_TEMPR21[62] ), .Y(
        OR2_41_Y));
    OR4 OR4_542 (.A(\R_DATA_TEMPR28[8] ), .B(\R_DATA_TEMPR29[8] ), .C(
        \R_DATA_TEMPR30[8] ), .D(\R_DATA_TEMPR31[8] ), .Y(OR4_542_Y));
    OR2 OR2_61 (.A(\R_DATA_TEMPR20[68] ), .B(\R_DATA_TEMPR21[68] ), .Y(
        OR2_61_Y));
    OR4 \OR4_R_DATA[4]  (.A(OR4_556_Y), .B(OR4_136_Y), .C(OR4_246_Y), 
        .D(OR4_312_Y), .Y(R_DATA[4]));
    OR4 OR4_135 (.A(\R_DATA_TEMPR12[41] ), .B(\R_DATA_TEMPR13[41] ), 
        .C(\R_DATA_TEMPR14[41] ), .D(\R_DATA_TEMPR15[41] ), .Y(
        OR4_135_Y));
    OR4 OR4_383 (.A(OR4_622_Y), .B(OR4_477_Y), .C(OR4_466_Y), .D(
        OR4_197_Y), .Y(OR4_383_Y));
    OR4 OR4_544 (.A(\R_DATA_TEMPR0[74] ), .B(\R_DATA_TEMPR1[74] ), .C(
        \R_DATA_TEMPR2[74] ), .D(\R_DATA_TEMPR3[74] ), .Y(OR4_544_Y));
    OR2 OR2_31 (.A(\R_DATA_TEMPR20[51] ), .B(\R_DATA_TEMPR21[51] ), .Y(
        OR2_31_Y));
    OR4 OR4_267 (.A(\R_DATA_TEMPR4[69] ), .B(\R_DATA_TEMPR5[69] ), .C(
        \R_DATA_TEMPR6[69] ), .D(\R_DATA_TEMPR7[69] ), .Y(OR4_267_Y));
    OR4 OR4_523 (.A(\R_DATA_TEMPR12[40] ), .B(\R_DATA_TEMPR13[40] ), 
        .C(\R_DATA_TEMPR14[40] ), .D(\R_DATA_TEMPR15[40] ), .Y(
        OR4_523_Y));
    OR4 OR4_437 (.A(OR4_128_Y), .B(OR2_35_Y), .C(\R_DATA_TEMPR22[22] ), 
        .D(\R_DATA_TEMPR23[22] ), .Y(OR4_437_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%7%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C1 (
        .A_DOUT({\R_DATA_TEMPR7[79] , \R_DATA_TEMPR7[78] , 
        \R_DATA_TEMPR7[77] , \R_DATA_TEMPR7[76] , \R_DATA_TEMPR7[75] , 
        \R_DATA_TEMPR7[74] , \R_DATA_TEMPR7[73] , \R_DATA_TEMPR7[72] , 
        \R_DATA_TEMPR7[71] , \R_DATA_TEMPR7[70] , \R_DATA_TEMPR7[69] , 
        \R_DATA_TEMPR7[68] , \R_DATA_TEMPR7[67] , \R_DATA_TEMPR7[66] , 
        \R_DATA_TEMPR7[65] , \R_DATA_TEMPR7[64] , \R_DATA_TEMPR7[63] , 
        \R_DATA_TEMPR7[62] , \R_DATA_TEMPR7[61] , \R_DATA_TEMPR7[60] })
        , .B_DOUT({\R_DATA_TEMPR7[59] , \R_DATA_TEMPR7[58] , 
        \R_DATA_TEMPR7[57] , \R_DATA_TEMPR7[56] , \R_DATA_TEMPR7[55] , 
        \R_DATA_TEMPR7[54] , \R_DATA_TEMPR7[53] , \R_DATA_TEMPR7[52] , 
        \R_DATA_TEMPR7[51] , \R_DATA_TEMPR7[50] , \R_DATA_TEMPR7[49] , 
        \R_DATA_TEMPR7[48] , \R_DATA_TEMPR7[47] , \R_DATA_TEMPR7[46] , 
        \R_DATA_TEMPR7[45] , \R_DATA_TEMPR7[44] , \R_DATA_TEMPR7[43] , 
        \R_DATA_TEMPR7[42] , \R_DATA_TEMPR7[41] , \R_DATA_TEMPR7[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[7][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[1] , 
        R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[1] , W_ADDR[10], W_ADDR[9]}), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_482 (.A(\R_DATA_TEMPR24[68] ), .B(\R_DATA_TEMPR25[68] ), 
        .C(\R_DATA_TEMPR26[68] ), .D(\R_DATA_TEMPR27[68] ), .Y(
        OR4_482_Y));
    OR4 OR4_167 (.A(\R_DATA_TEMPR8[17] ), .B(\R_DATA_TEMPR9[17] ), .C(
        \R_DATA_TEMPR10[17] ), .D(\R_DATA_TEMPR11[17] ), .Y(OR4_167_Y));
    OR4 OR4_705 (.A(OR4_146_Y), .B(OR2_43_Y), .C(\R_DATA_TEMPR22[76] ), 
        .D(\R_DATA_TEMPR23[76] ), .Y(OR4_705_Y));
    OR4 OR4_607 (.A(OR4_177_Y), .B(OR4_410_Y), .C(OR4_719_Y), .D(
        OR4_296_Y), .Y(OR4_607_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%21%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C1 (
        .A_DOUT({\R_DATA_TEMPR21[79] , \R_DATA_TEMPR21[78] , 
        \R_DATA_TEMPR21[77] , \R_DATA_TEMPR21[76] , 
        \R_DATA_TEMPR21[75] , \R_DATA_TEMPR21[74] , 
        \R_DATA_TEMPR21[73] , \R_DATA_TEMPR21[72] , 
        \R_DATA_TEMPR21[71] , \R_DATA_TEMPR21[70] , 
        \R_DATA_TEMPR21[69] , \R_DATA_TEMPR21[68] , 
        \R_DATA_TEMPR21[67] , \R_DATA_TEMPR21[66] , 
        \R_DATA_TEMPR21[65] , \R_DATA_TEMPR21[64] , 
        \R_DATA_TEMPR21[63] , \R_DATA_TEMPR21[62] , 
        \R_DATA_TEMPR21[61] , \R_DATA_TEMPR21[60] }), .B_DOUT({
        \R_DATA_TEMPR21[59] , \R_DATA_TEMPR21[58] , 
        \R_DATA_TEMPR21[57] , \R_DATA_TEMPR21[56] , 
        \R_DATA_TEMPR21[55] , \R_DATA_TEMPR21[54] , 
        \R_DATA_TEMPR21[53] , \R_DATA_TEMPR21[52] , 
        \R_DATA_TEMPR21[51] , \R_DATA_TEMPR21[50] , 
        \R_DATA_TEMPR21[49] , \R_DATA_TEMPR21[48] , 
        \R_DATA_TEMPR21[47] , \R_DATA_TEMPR21[46] , 
        \R_DATA_TEMPR21[45] , \R_DATA_TEMPR21[44] , 
        \R_DATA_TEMPR21[43] , \R_DATA_TEMPR21[42] , 
        \R_DATA_TEMPR21[41] , \R_DATA_TEMPR21[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[21][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_489 (.A(\R_DATA_TEMPR12[77] ), .B(\R_DATA_TEMPR13[77] ), 
        .C(\R_DATA_TEMPR14[77] ), .D(\R_DATA_TEMPR15[77] ), .Y(
        OR4_489_Y));
    OR4 OR4_706 (.A(\R_DATA_TEMPR24[11] ), .B(\R_DATA_TEMPR25[11] ), 
        .C(\R_DATA_TEMPR26[11] ), .D(\R_DATA_TEMPR27[11] ), .Y(
        OR4_706_Y));
    OR4 OR4_186 (.A(\R_DATA_TEMPR24[67] ), .B(\R_DATA_TEMPR25[67] ), 
        .C(\R_DATA_TEMPR26[67] ), .D(\R_DATA_TEMPR27[67] ), .Y(
        OR4_186_Y));
    OR4 OR4_677 (.A(OR4_427_Y), .B(OR2_68_Y), .C(\R_DATA_TEMPR22[1] ), 
        .D(\R_DATA_TEMPR23[1] ), .Y(OR4_677_Y));
    OR4 OR4_235 (.A(OR4_89_Y), .B(OR2_57_Y), .C(\R_DATA_TEMPR22[73] ), 
        .D(\R_DATA_TEMPR23[73] ), .Y(OR4_235_Y));
    OR4 OR4_341 (.A(OR4_559_Y), .B(OR2_22_Y), .C(\R_DATA_TEMPR22[41] ), 
        .D(\R_DATA_TEMPR23[41] ), .Y(OR4_341_Y));
    OR2 OR2_29 (.A(\R_DATA_TEMPR20[18] ), .B(\R_DATA_TEMPR21[18] ), .Y(
        OR2_29_Y));
    OR4 OR4_264 (.A(\R_DATA_TEMPR28[30] ), .B(\R_DATA_TEMPR29[30] ), 
        .C(\R_DATA_TEMPR30[30] ), .D(\R_DATA_TEMPR31[30] ), .Y(
        OR4_264_Y));
    OR4 OR4_656 (.A(\R_DATA_TEMPR0[12] ), .B(\R_DATA_TEMPR1[12] ), .C(
        \R_DATA_TEMPR2[12] ), .D(\R_DATA_TEMPR3[12] ), .Y(OR4_656_Y));
    OR4 OR4_440 (.A(OR4_41_Y), .B(OR2_48_Y), .C(\R_DATA_TEMPR22[49] ), 
        .D(\R_DATA_TEMPR23[49] ), .Y(OR4_440_Y));
    OR4 OR4_293 (.A(\R_DATA_TEMPR16[3] ), .B(\R_DATA_TEMPR17[3] ), .C(
        \R_DATA_TEMPR18[3] ), .D(\R_DATA_TEMPR19[3] ), .Y(OR4_293_Y));
    OR4 OR4_388 (.A(\R_DATA_TEMPR28[66] ), .B(\R_DATA_TEMPR29[66] ), 
        .C(\R_DATA_TEMPR30[66] ), .D(\R_DATA_TEMPR31[66] ), .Y(
        OR4_388_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%13%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0 (
        .A_DOUT({\R_DATA_TEMPR13[39] , \R_DATA_TEMPR13[38] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR13[36] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR13[34] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR13[32] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR13[30] , 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR13[28] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR13[26] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR13[24] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR13[22] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR13[20] }), .B_DOUT({
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR13[18] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR13[16] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR13[14] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR13[12] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR13[10] , 
        \R_DATA_TEMPR13[9] , \R_DATA_TEMPR13[8] , \R_DATA_TEMPR13[7] , 
        \R_DATA_TEMPR13[6] , \R_DATA_TEMPR13[5] , \R_DATA_TEMPR13[4] , 
        \R_DATA_TEMPR13[3] , \R_DATA_TEMPR13[2] , \R_DATA_TEMPR13[1] , 
        \R_DATA_TEMPR13[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_115 (.A(OR4_404_Y), .B(OR4_94_Y), .C(OR4_127_Y), .D(
        OR4_503_Y), .Y(OR4_115_Y));
    OR4 OR4_66 (.A(OR4_386_Y), .B(OR2_55_Y), .C(\R_DATA_TEMPR22[19] ), 
        .D(\R_DATA_TEMPR23[19] ), .Y(OR4_66_Y));
    OR4 OR4_433 (.A(OR4_331_Y), .B(OR2_71_Y), .C(\R_DATA_TEMPR22[27] ), 
        .D(\R_DATA_TEMPR23[27] ), .Y(OR4_433_Y));
    OR4 OR4_417 (.A(\R_DATA_TEMPR24[9] ), .B(\R_DATA_TEMPR25[9] ), .C(
        \R_DATA_TEMPR26[9] ), .D(\R_DATA_TEMPR27[9] ), .Y(OR4_417_Y));
    OR4 OR4_631 (.A(\R_DATA_TEMPR16[14] ), .B(\R_DATA_TEMPR17[14] ), 
        .C(\R_DATA_TEMPR18[14] ), .D(\R_DATA_TEMPR19[14] ), .Y(
        OR4_631_Y));
    CFG2 #( .INIT(4'h1) )  CFG2_4 (.A(W_ADDR[12]), .B(W_ADDR[11]), .Y(
        CFG2_4_Y));
    OR4 OR4_365 (.A(\R_DATA_TEMPR8[38] ), .B(\R_DATA_TEMPR9[38] ), .C(
        \R_DATA_TEMPR10[38] ), .D(\R_DATA_TEMPR11[38] ), .Y(OR4_365_Y));
    OR4 OR4_238 (.A(\R_DATA_TEMPR0[53] ), .B(\R_DATA_TEMPR1[53] ), .C(
        \R_DATA_TEMPR2[53] ), .D(\R_DATA_TEMPR3[53] ), .Y(OR4_238_Y));
    OR2 OR2_8 (.A(\R_DATA_TEMPR20[45] ), .B(\R_DATA_TEMPR21[45] ), .Y(
        OR2_8_Y));
    OR4 \OR4_R_DATA[52]  (.A(OR4_62_Y), .B(OR4_44_Y), .C(OR4_671_Y), 
        .D(OR4_344_Y), .Y(R_DATA[52]));
    OR4 OR4_189 (.A(OR4_59_Y), .B(OR4_226_Y), .C(OR4_295_Y), .D(
        OR4_93_Y), .Y(OR4_189_Y));
    OR4 OR4_0 (.A(\R_DATA_TEMPR8[62] ), .B(\R_DATA_TEMPR9[62] ), .C(
        \R_DATA_TEMPR10[62] ), .D(\R_DATA_TEMPR11[62] ), .Y(OR4_0_Y));
    OR4 OR4_207 (.A(\R_DATA_TEMPR8[40] ), .B(\R_DATA_TEMPR9[40] ), .C(
        \R_DATA_TEMPR10[40] ), .D(\R_DATA_TEMPR11[40] ), .Y(OR4_207_Y));
    OR4 OR4_215 (.A(\R_DATA_TEMPR12[2] ), .B(\R_DATA_TEMPR13[2] ), .C(
        \R_DATA_TEMPR14[2] ), .D(\R_DATA_TEMPR15[2] ), .Y(OR4_215_Y));
    OR4 OR4_107 (.A(OR4_321_Y), .B(OR4_575_Y), .C(OR4_516_Y), .D(
        OR4_228_Y), .Y(OR4_107_Y));
    OR4 OR4_277 (.A(OR4_517_Y), .B(OR4_643_Y), .C(OR4_640_Y), .D(
        OR4_33_Y), .Y(OR4_277_Y));
    OR4 OR4_698 (.A(OR4_74_Y), .B(OR2_40_Y), .C(\R_DATA_TEMPR22[20] ), 
        .D(\R_DATA_TEMPR23[20] ), .Y(OR4_698_Y));
    OR4 OR4_95 (.A(\R_DATA_TEMPR4[67] ), .B(\R_DATA_TEMPR5[67] ), .C(
        \R_DATA_TEMPR6[67] ), .D(\R_DATA_TEMPR7[67] ), .Y(OR4_95_Y));
    OR2 OR2_22 (.A(\R_DATA_TEMPR20[41] ), .B(\R_DATA_TEMPR21[41] ), .Y(
        OR2_22_Y));
    OR4 OR4_177 (.A(\R_DATA_TEMPR0[49] ), .B(\R_DATA_TEMPR1[49] ), .C(
        \R_DATA_TEMPR2[49] ), .D(\R_DATA_TEMPR3[49] ), .Y(OR4_177_Y));
    OR2 OR2_79 (.A(\R_DATA_TEMPR20[29] ), .B(\R_DATA_TEMPR21[29] ), .Y(
        OR2_79_Y));
    OR4 \OR4_R_DATA[34]  (.A(OR4_122_Y), .B(OR4_604_Y), .C(OR4_243_Y), 
        .D(OR4_547_Y), .Y(R_DATA[34]));
    OR4 OR4_349 (.A(\R_DATA_TEMPR28[50] ), .B(\R_DATA_TEMPR29[50] ), 
        .C(\R_DATA_TEMPR30[50] ), .D(\R_DATA_TEMPR31[50] ), .Y(
        OR4_349_Y));
    OR4 OR4_692 (.A(\R_DATA_TEMPR28[27] ), .B(\R_DATA_TEMPR29[27] ), 
        .C(\R_DATA_TEMPR30[27] ), .D(\R_DATA_TEMPR31[27] ), .Y(
        OR4_692_Y));
    OR4 OR4_703 (.A(\R_DATA_TEMPR0[30] ), .B(\R_DATA_TEMPR1[30] ), .C(
        \R_DATA_TEMPR2[30] ), .D(\R_DATA_TEMPR3[30] ), .Y(OR4_703_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%10%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C1 (
        .A_DOUT({\R_DATA_TEMPR10[79] , \R_DATA_TEMPR10[78] , 
        \R_DATA_TEMPR10[77] , \R_DATA_TEMPR10[76] , 
        \R_DATA_TEMPR10[75] , \R_DATA_TEMPR10[74] , 
        \R_DATA_TEMPR10[73] , \R_DATA_TEMPR10[72] , 
        \R_DATA_TEMPR10[71] , \R_DATA_TEMPR10[70] , 
        \R_DATA_TEMPR10[69] , \R_DATA_TEMPR10[68] , 
        \R_DATA_TEMPR10[67] , \R_DATA_TEMPR10[66] , 
        \R_DATA_TEMPR10[65] , \R_DATA_TEMPR10[64] , 
        \R_DATA_TEMPR10[63] , \R_DATA_TEMPR10[62] , 
        \R_DATA_TEMPR10[61] , \R_DATA_TEMPR10[60] }), .B_DOUT({
        \R_DATA_TEMPR10[59] , \R_DATA_TEMPR10[58] , 
        \R_DATA_TEMPR10[57] , \R_DATA_TEMPR10[56] , 
        \R_DATA_TEMPR10[55] , \R_DATA_TEMPR10[54] , 
        \R_DATA_TEMPR10[53] , \R_DATA_TEMPR10[52] , 
        \R_DATA_TEMPR10[51] , \R_DATA_TEMPR10[50] , 
        \R_DATA_TEMPR10[49] , \R_DATA_TEMPR10[48] , 
        \R_DATA_TEMPR10[47] , \R_DATA_TEMPR10[46] , 
        \R_DATA_TEMPR10[45] , \R_DATA_TEMPR10[44] , 
        \R_DATA_TEMPR10[43] , \R_DATA_TEMPR10[42] , 
        \R_DATA_TEMPR10[41] , \R_DATA_TEMPR10[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[10][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_223 (.A(\R_DATA_TEMPR0[17] ), .B(\R_DATA_TEMPR1[17] ), .C(
        \R_DATA_TEMPR2[17] ), .D(\R_DATA_TEMPR3[17] ), .Y(OR4_223_Y));
    OR4 OR4_204 (.A(\R_DATA_TEMPR0[15] ), .B(\R_DATA_TEMPR1[15] ), .C(
        \R_DATA_TEMPR2[15] ), .D(\R_DATA_TEMPR3[15] ), .Y(OR4_204_Y));
    OR4 OR4_354 (.A(\R_DATA_TEMPR0[35] ), .B(\R_DATA_TEMPR1[35] ), .C(
        \R_DATA_TEMPR2[35] ), .D(\R_DATA_TEMPR3[35] ), .Y(OR4_354_Y));
    OR2 OR2_19 (.A(\R_DATA_TEMPR20[6] ), .B(\R_DATA_TEMPR21[6] ), .Y(
        OR2_19_Y));
    OR4 OR4_665 (.A(\R_DATA_TEMPR0[1] ), .B(\R_DATA_TEMPR1[1] ), .C(
        \R_DATA_TEMPR2[1] ), .D(\R_DATA_TEMPR3[1] ), .Y(OR4_665_Y));
    OR4 OR4_413 (.A(\R_DATA_TEMPR8[68] ), .B(\R_DATA_TEMPR9[68] ), .C(
        \R_DATA_TEMPR10[68] ), .D(\R_DATA_TEMPR11[68] ), .Y(OR4_413_Y));
    OR4 OR4_611 (.A(OR4_116_Y), .B(OR4_709_Y), .C(OR4_693_Y), .D(
        OR4_409_Y), .Y(OR4_611_Y));
    OR4 OR4_151 (.A(\R_DATA_TEMPR0[27] ), .B(\R_DATA_TEMPR1[27] ), .C(
        \R_DATA_TEMPR2[27] ), .D(\R_DATA_TEMPR3[27] ), .Y(OR4_151_Y));
    OR4 OR4_274 (.A(\R_DATA_TEMPR28[25] ), .B(\R_DATA_TEMPR29[25] ), 
        .C(\R_DATA_TEMPR30[25] ), .D(\R_DATA_TEMPR31[25] ), .Y(
        OR4_274_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%31%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0 (
        .A_DOUT({\R_DATA_TEMPR31[39] , \R_DATA_TEMPR31[38] , 
        \R_DATA_TEMPR31[37] , \R_DATA_TEMPR31[36] , 
        \R_DATA_TEMPR31[35] , \R_DATA_TEMPR31[34] , 
        \R_DATA_TEMPR31[33] , \R_DATA_TEMPR31[32] , 
        \R_DATA_TEMPR31[31] , \R_DATA_TEMPR31[30] , 
        \R_DATA_TEMPR31[29] , \R_DATA_TEMPR31[28] , 
        \R_DATA_TEMPR31[27] , \R_DATA_TEMPR31[26] , 
        \R_DATA_TEMPR31[25] , \R_DATA_TEMPR31[24] , 
        \R_DATA_TEMPR31[23] , \R_DATA_TEMPR31[22] , 
        \R_DATA_TEMPR31[21] , \R_DATA_TEMPR31[20] }), .B_DOUT({
        \R_DATA_TEMPR31[19] , \R_DATA_TEMPR31[18] , 
        \R_DATA_TEMPR31[17] , \R_DATA_TEMPR31[16] , 
        \R_DATA_TEMPR31[15] , \R_DATA_TEMPR31[14] , 
        \R_DATA_TEMPR31[13] , \R_DATA_TEMPR31[12] , 
        \R_DATA_TEMPR31[11] , \R_DATA_TEMPR31[10] , 
        \R_DATA_TEMPR31[9] , \R_DATA_TEMPR31[8] , \R_DATA_TEMPR31[7] , 
        \R_DATA_TEMPR31[6] , \R_DATA_TEMPR31[5] , \R_DATA_TEMPR31[4] , 
        \R_DATA_TEMPR31[3] , \R_DATA_TEMPR31[2] , \R_DATA_TEMPR31[1] , 
        \R_DATA_TEMPR31[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_218 (.A(OR4_492_Y), .B(OR4_7_Y), .C(OR4_318_Y), .D(
        OR4_617_Y), .Y(OR4_218_Y));
    OR4 \OR4_R_DATA[22]  (.A(OR4_462_Y), .B(OR4_437_Y), .C(OR4_339_Y), 
        .D(OR4_18_Y), .Y(R_DATA[22]));
    OR4 \OR4_R_DATA[53]  (.A(OR4_712_Y), .B(OR4_521_Y), .C(OR4_493_Y), 
        .D(OR4_470_Y), .Y(R_DATA[53]));
    OR4 OR4_60 (.A(\R_DATA_TEMPR24[14] ), .B(\R_DATA_TEMPR25[14] ), .C(
        \R_DATA_TEMPR26[14] ), .D(\R_DATA_TEMPR27[14] ), .Y(OR4_60_Y));
    OR4 OR4_531 (.A(\R_DATA_TEMPR28[38] ), .B(\R_DATA_TEMPR29[38] ), 
        .C(\R_DATA_TEMPR30[38] ), .D(\R_DATA_TEMPR31[38] ), .Y(
        OR4_531_Y));
    OR4 OR4_67 (.A(OR4_354_Y), .B(OR4_50_Y), .C(OR4_77_Y), .D(
        OR4_449_Y), .Y(OR4_67_Y));
    OR4 OR4_687 (.A(\R_DATA_TEMPR4[66] ), .B(\R_DATA_TEMPR5[66] ), .C(
        \R_DATA_TEMPR6[66] ), .D(\R_DATA_TEMPR7[66] ), .Y(OR4_687_Y));
    OR4 OR4_305 (.A(\R_DATA_TEMPR0[42] ), .B(\R_DATA_TEMPR1[42] ), .C(
        \R_DATA_TEMPR2[42] ), .D(\R_DATA_TEMPR3[42] ), .Y(OR4_305_Y));
    OR4 OR4_451 (.A(\R_DATA_TEMPR8[44] ), .B(\R_DATA_TEMPR9[44] ), .C(
        \R_DATA_TEMPR10[44] ), .D(\R_DATA_TEMPR11[44] ), .Y(OR4_451_Y));
    OR4 OR4_458 (.A(\R_DATA_TEMPR0[29] ), .B(\R_DATA_TEMPR1[29] ), .C(
        \R_DATA_TEMPR2[29] ), .D(\R_DATA_TEMPR3[29] ), .Y(OR4_458_Y));
    OR4 OR4_628 (.A(OR4_496_Y), .B(OR2_70_Y), .C(\R_DATA_TEMPR22[43] ), 
        .D(\R_DATA_TEMPR23[43] ), .Y(OR4_628_Y));
    OR4 OR4_375 (.A(\R_DATA_TEMPR16[9] ), .B(\R_DATA_TEMPR17[9] ), .C(
        \R_DATA_TEMPR18[9] ), .D(\R_DATA_TEMPR19[9] ), .Y(OR4_375_Y));
    OR2 OR2_72 (.A(\R_DATA_TEMPR20[70] ), .B(\R_DATA_TEMPR21[70] ), .Y(
        OR2_72_Y));
    OR4 OR4_660 (.A(OR4_544_Y), .B(OR4_699_Y), .C(OR4_48_Y), .D(
        OR4_581_Y), .Y(OR4_660_Y));
    OR4 OR4_622 (.A(\R_DATA_TEMPR0[23] ), .B(\R_DATA_TEMPR1[23] ), .C(
        \R_DATA_TEMPR2[23] ), .D(\R_DATA_TEMPR3[23] ), .Y(OR4_622_Y));
    OR4 OR4_232 (.A(\R_DATA_TEMPR0[44] ), .B(\R_DATA_TEMPR1[44] ), .C(
        \R_DATA_TEMPR2[44] ), .D(\R_DATA_TEMPR3[44] ), .Y(OR4_232_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[4]  (.A(CFG2_3_Y), .B(
        R_ADDR[13]), .C(R_EN), .Y(\BLKY2[4] ));
    OR4 \OR4_R_DATA[15]  (.A(OR4_636_Y), .B(OR4_265_Y), .C(OR4_535_Y), 
        .D(OR4_320_Y), .Y(R_DATA[15]));
    OR4 OR4_543 (.A(\R_DATA_TEMPR8[10] ), .B(\R_DATA_TEMPR9[10] ), .C(
        \R_DATA_TEMPR10[10] ), .D(\R_DATA_TEMPR11[10] ), .Y(OR4_543_Y));
    OR4 OR4_45 (.A(\R_DATA_TEMPR28[72] ), .B(\R_DATA_TEMPR29[72] ), .C(
        \R_DATA_TEMPR30[72] ), .D(\R_DATA_TEMPR31[72] ), .Y(OR4_45_Y));
    OR4 OR4_367 (.A(\R_DATA_TEMPR8[11] ), .B(\R_DATA_TEMPR9[11] ), .C(
        \R_DATA_TEMPR10[11] ), .D(\R_DATA_TEMPR11[11] ), .Y(OR4_367_Y));
    OR4 OR4_160 (.A(\R_DATA_TEMPR8[46] ), .B(\R_DATA_TEMPR9[46] ), .C(
        \R_DATA_TEMPR10[46] ), .D(\R_DATA_TEMPR11[46] ), .Y(OR4_160_Y));
    OR2 OR2_12 (.A(\R_DATA_TEMPR20[10] ), .B(\R_DATA_TEMPR21[10] ), .Y(
        OR2_12_Y));
    OR4 OR4_702 (.A(\R_DATA_TEMPR12[0] ), .B(\R_DATA_TEMPR13[0] ), .C(
        \R_DATA_TEMPR14[0] ), .D(\R_DATA_TEMPR15[0] ), .Y(OR4_702_Y));
    OR4 OR4_559 (.A(\R_DATA_TEMPR16[41] ), .B(\R_DATA_TEMPR17[41] ), 
        .C(\R_DATA_TEMPR18[41] ), .D(\R_DATA_TEMPR19[41] ), .Y(
        OR4_559_Y));
    OR4 OR4_550 (.A(\R_DATA_TEMPR12[24] ), .B(\R_DATA_TEMPR13[24] ), 
        .C(\R_DATA_TEMPR14[24] ), .D(\R_DATA_TEMPR15[24] ), .Y(
        OR4_550_Y));
    OR4 \OR4_R_DATA[23]  (.A(OR4_383_Y), .B(OR4_206_Y), .C(OR4_164_Y), 
        .D(OR4_139_Y), .Y(R_DATA[23]));
    OR4 OR4_330 (.A(OR4_684_Y), .B(OR4_471_Y), .C(OR4_509_Y), .D(
        OR4_645_Y), .Y(OR4_330_Y));
    OR4 OR4_605 (.A(OR4_161_Y), .B(OR4_583_Y), .C(OR4_615_Y), .D(
        OR4_269_Y), .Y(OR4_605_Y));
    OR4 OR4_511 (.A(\R_DATA_TEMPR0[24] ), .B(\R_DATA_TEMPR1[24] ), .C(
        \R_DATA_TEMPR2[24] ), .D(\R_DATA_TEMPR3[24] ), .Y(OR4_511_Y));
    OR4 OR4_696 (.A(\R_DATA_TEMPR0[7] ), .B(\R_DATA_TEMPR1[7] ), .C(
        \R_DATA_TEMPR2[7] ), .D(\R_DATA_TEMPR3[7] ), .Y(OR4_696_Y));
    OR4 OR4_675 (.A(\R_DATA_TEMPR8[32] ), .B(\R_DATA_TEMPR9[32] ), .C(
        \R_DATA_TEMPR10[32] ), .D(\R_DATA_TEMPR11[32] ), .Y(OR4_675_Y));
    OR4 OR4_287 (.A(\R_DATA_TEMPR12[46] ), .B(\R_DATA_TEMPR13[46] ), 
        .C(\R_DATA_TEMPR14[46] ), .D(\R_DATA_TEMPR15[46] ), .Y(
        OR4_287_Y));
    OR4 OR4_86 (.A(\R_DATA_TEMPR8[4] ), .B(\R_DATA_TEMPR9[4] ), .C(
        \R_DATA_TEMPR10[4] ), .D(\R_DATA_TEMPR11[4] ), .Y(OR4_86_Y));
    OR4 OR4_33 (.A(\R_DATA_TEMPR12[51] ), .B(\R_DATA_TEMPR13[51] ), .C(
        \R_DATA_TEMPR14[51] ), .D(\R_DATA_TEMPR15[51] ), .Y(OR4_33_Y));
    OR4 OR4_168 (.A(OR4_92_Y), .B(OR4_327_Y), .C(OR4_179_Y), .D(
        OR4_174_Y), .Y(OR4_168_Y));
    OR4 OR4_187 (.A(\R_DATA_TEMPR16[11] ), .B(\R_DATA_TEMPR17[11] ), 
        .C(\R_DATA_TEMPR18[11] ), .D(\R_DATA_TEMPR19[11] ), .Y(
        OR4_187_Y));
    OR2 OR2_46 (.A(\R_DATA_TEMPR20[2] ), .B(\R_DATA_TEMPR21[2] ), .Y(
        OR2_46_Y));
    OR4 OR4_212 (.A(\R_DATA_TEMPR8[18] ), .B(\R_DATA_TEMPR9[18] ), .C(
        \R_DATA_TEMPR10[18] ), .D(\R_DATA_TEMPR11[18] ), .Y(OR4_212_Y));
    OR4 OR4_353 (.A(\R_DATA_TEMPR28[7] ), .B(\R_DATA_TEMPR29[7] ), .C(
        \R_DATA_TEMPR30[7] ), .D(\R_DATA_TEMPR31[7] ), .Y(OR4_353_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%6%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0 (
        .A_DOUT({\R_DATA_TEMPR6[39] , \R_DATA_TEMPR6[38] , 
        \R_DATA_TEMPR6[37] , \R_DATA_TEMPR6[36] , \R_DATA_TEMPR6[35] , 
        \R_DATA_TEMPR6[34] , \R_DATA_TEMPR6[33] , \R_DATA_TEMPR6[32] , 
        \R_DATA_TEMPR6[31] , \R_DATA_TEMPR6[30] , \R_DATA_TEMPR6[29] , 
        \R_DATA_TEMPR6[28] , \R_DATA_TEMPR6[27] , \R_DATA_TEMPR6[26] , 
        \R_DATA_TEMPR6[25] , \R_DATA_TEMPR6[24] , \R_DATA_TEMPR6[23] , 
        \R_DATA_TEMPR6[22] , \R_DATA_TEMPR6[21] , \R_DATA_TEMPR6[20] })
        , .B_DOUT({\R_DATA_TEMPR6[19] , \R_DATA_TEMPR6[18] , 
        \R_DATA_TEMPR6[17] , \R_DATA_TEMPR6[16] , \R_DATA_TEMPR6[15] , 
        \R_DATA_TEMPR6[14] , \R_DATA_TEMPR6[13] , \R_DATA_TEMPR6[12] , 
        \R_DATA_TEMPR6[11] , \R_DATA_TEMPR6[10] , \R_DATA_TEMPR6[9] , 
        \R_DATA_TEMPR6[8] , \R_DATA_TEMPR6[7] , \R_DATA_TEMPR6[6] , 
        \R_DATA_TEMPR6[5] , \R_DATA_TEMPR6[4] , \R_DATA_TEMPR6[3] , 
        \R_DATA_TEMPR6[2] , \R_DATA_TEMPR6[1] , \R_DATA_TEMPR6[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[6][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[45]  (.A(OR4_282_Y), .B(OR4_627_Y), .C(OR4_194_Y), 
        .D(OR4_707_Y), .Y(R_DATA[45]));
    OR4 OR4_600 (.A(\R_DATA_TEMPR4[60] ), .B(\R_DATA_TEMPR5[60] ), .C(
        \R_DATA_TEMPR6[60] ), .D(\R_DATA_TEMPR7[60] ), .Y(OR4_600_Y));
    OR4 OR4_452 (.A(\R_DATA_TEMPR24[0] ), .B(\R_DATA_TEMPR25[0] ), .C(
        \R_DATA_TEMPR26[0] ), .D(\R_DATA_TEMPR27[0] ), .Y(OR4_452_Y));
    OR4 OR4_284 (.A(\R_DATA_TEMPR12[15] ), .B(\R_DATA_TEMPR13[15] ), 
        .C(\R_DATA_TEMPR14[15] ), .D(\R_DATA_TEMPR15[15] ), .Y(
        OR4_284_Y));
    OR4 OR4_310 (.A(\R_DATA_TEMPR12[32] ), .B(\R_DATA_TEMPR13[32] ), 
        .C(\R_DATA_TEMPR14[32] ), .D(\R_DATA_TEMPR15[32] ), .Y(
        OR4_310_Y));
    OR4 OR4_5 (.A(\R_DATA_TEMPR12[67] ), .B(\R_DATA_TEMPR13[67] ), .C(
        \R_DATA_TEMPR14[67] ), .D(\R_DATA_TEMPR15[67] ), .Y(OR4_5_Y));
    OR4 OR4_670 (.A(OR4_563_Y), .B(OR2_58_Y), .C(\R_DATA_TEMPR22[37] ), 
        .D(\R_DATA_TEMPR23[37] ), .Y(OR4_670_Y));
    OR2 OR2_66 (.A(\R_DATA_TEMPR20[56] ), .B(\R_DATA_TEMPR21[56] ), .Y(
        OR2_66_Y));
    OR4 OR4_459 (.A(\R_DATA_TEMPR24[7] ), .B(\R_DATA_TEMPR25[7] ), .C(
        \R_DATA_TEMPR26[7] ), .D(\R_DATA_TEMPR27[7] ), .Y(OR4_459_Y));
    OR4 OR4_307 (.A(\R_DATA_TEMPR8[21] ), .B(\R_DATA_TEMPR9[21] ), .C(
        \R_DATA_TEMPR10[21] ), .D(\R_DATA_TEMPR11[21] ), .Y(OR4_307_Y));
    OR4 OR4_100 (.A(\R_DATA_TEMPR0[8] ), .B(\R_DATA_TEMPR1[8] ), .C(
        \R_DATA_TEMPR2[8] ), .D(\R_DATA_TEMPR3[8] ), .Y(OR4_100_Y));
    OR4 OR4_99 (.A(\R_DATA_TEMPR16[0] ), .B(\R_DATA_TEMPR17[0] ), .C(
        \R_DATA_TEMPR18[0] ), .D(\R_DATA_TEMPR19[0] ), .Y(OR4_99_Y));
    OR4 OR4_156 (.A(OR4_570_Y), .B(OR2_77_Y), .C(\R_DATA_TEMPR22[42] ), 
        .D(\R_DATA_TEMPR23[42] ), .Y(OR4_156_Y));
    OR4 OR4_535 (.A(\R_DATA_TEMPR24[15] ), .B(\R_DATA_TEMPR25[15] ), 
        .C(\R_DATA_TEMPR26[15] ), .D(\R_DATA_TEMPR27[15] ), .Y(
        OR4_535_Y));
    OR2 OR2_36 (.A(\R_DATA_TEMPR20[34] ), .B(\R_DATA_TEMPR21[34] ), .Y(
        OR2_36_Y));
    OR4 OR4_68 (.A(\R_DATA_TEMPR24[26] ), .B(\R_DATA_TEMPR25[26] ), .C(
        \R_DATA_TEMPR26[26] ), .D(\R_DATA_TEMPR27[26] ), .Y(OR4_68_Y));
    OR2 OR2_24 (.A(\R_DATA_TEMPR20[23] ), .B(\R_DATA_TEMPR21[23] ), .Y(
        OR2_24_Y));
    OR4 OR4_377 (.A(\R_DATA_TEMPR16[38] ), .B(\R_DATA_TEMPR17[38] ), 
        .C(\R_DATA_TEMPR18[38] ), .D(\R_DATA_TEMPR19[38] ), .Y(
        OR4_377_Y));
    OR4 OR4_170 (.A(OR4_415_Y), .B(OR4_540_Y), .C(OR4_538_Y), .D(
        OR4_653_Y), .Y(OR4_170_Y));
    OR4 OR4_708 (.A(OR4_175_Y), .B(OR2_26_Y), .C(\R_DATA_TEMPR22[54] ), 
        .D(\R_DATA_TEMPR23[54] ), .Y(OR4_708_Y));
    OR4 OR4_626 (.A(\R_DATA_TEMPR0[72] ), .B(\R_DATA_TEMPR1[72] ), .C(
        \R_DATA_TEMPR2[72] ), .D(\R_DATA_TEMPR3[72] ), .Y(OR4_626_Y));
    OR4 OR4_31 (.A(\R_DATA_TEMPR4[63] ), .B(\R_DATA_TEMPR5[63] ), .C(
        \R_DATA_TEMPR6[63] ), .D(\R_DATA_TEMPR7[63] ), .Y(OR4_31_Y));
    OR4 \OR4_R_DATA[65]  (.A(OR4_115_Y), .B(OR4_468_Y), .C(OR4_28_Y), 
        .D(OR4_546_Y), .Y(R_DATA[65]));
    OR4 OR4_633 (.A(OR4_405_Y), .B(OR4_268_Y), .C(OR4_132_Y), .D(
        OR4_172_Y), .Y(OR4_633_Y));
    OR4 \OR4_R_DATA[31]  (.A(OR4_170_Y), .B(OR4_126_Y), .C(OR4_142_Y), 
        .D(OR4_648_Y), .Y(R_DATA[31]));
    OR4 OR4_385 (.A(\R_DATA_TEMPR8[67] ), .B(\R_DATA_TEMPR9[67] ), .C(
        \R_DATA_TEMPR10[67] ), .D(\R_DATA_TEMPR11[67] ), .Y(OR4_385_Y));
    OR4 OR4_243 (.A(\R_DATA_TEMPR24[34] ), .B(\R_DATA_TEMPR25[34] ), 
        .C(\R_DATA_TEMPR26[34] ), .D(\R_DATA_TEMPR27[34] ), .Y(
        OR4_243_Y));
    OR4 OR4_394 (.A(\R_DATA_TEMPR16[61] ), .B(\R_DATA_TEMPR17[61] ), 
        .C(\R_DATA_TEMPR18[61] ), .D(\R_DATA_TEMPR19[61] ), .Y(
        OR4_394_Y));
    OR4 OR4_358 (.A(OR4_490_Y), .B(OR2_46_Y), .C(\R_DATA_TEMPR22[2] ), 
        .D(\R_DATA_TEMPR23[2] ), .Y(OR4_358_Y));
    OR4 OR4_80 (.A(\R_DATA_TEMPR12[22] ), .B(\R_DATA_TEMPR13[22] ), .C(
        \R_DATA_TEMPR14[22] ), .D(\R_DATA_TEMPR15[22] ), .Y(OR4_80_Y));
    OR4 OR4_108 (.A(\R_DATA_TEMPR12[72] ), .B(\R_DATA_TEMPR13[72] ), 
        .C(\R_DATA_TEMPR14[72] ), .D(\R_DATA_TEMPR15[72] ), .Y(
        OR4_108_Y));
    OR4 OR4_191 (.A(OR4_683_Y), .B(OR4_537_Y), .C(OR4_413_Y), .D(
        OR4_444_Y), .Y(OR4_191_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%12%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C1 (
        .A_DOUT({\R_DATA_TEMPR12[79] , \R_DATA_TEMPR12[78] , 
        \R_DATA_TEMPR12[77] , \R_DATA_TEMPR12[76] , 
        \R_DATA_TEMPR12[75] , \R_DATA_TEMPR12[74] , 
        \R_DATA_TEMPR12[73] , \R_DATA_TEMPR12[72] , 
        \R_DATA_TEMPR12[71] , \R_DATA_TEMPR12[70] , 
        \R_DATA_TEMPR12[69] , \R_DATA_TEMPR12[68] , 
        \R_DATA_TEMPR12[67] , \R_DATA_TEMPR12[66] , 
        \R_DATA_TEMPR12[65] , \R_DATA_TEMPR12[64] , 
        \R_DATA_TEMPR12[63] , \R_DATA_TEMPR12[62] , 
        \R_DATA_TEMPR12[61] , \R_DATA_TEMPR12[60] }), .B_DOUT({
        \R_DATA_TEMPR12[59] , \R_DATA_TEMPR12[58] , 
        \R_DATA_TEMPR12[57] , \R_DATA_TEMPR12[56] , 
        \R_DATA_TEMPR12[55] , \R_DATA_TEMPR12[54] , 
        \R_DATA_TEMPR12[53] , \R_DATA_TEMPR12[52] , 
        \R_DATA_TEMPR12[51] , \R_DATA_TEMPR12[50] , 
        \R_DATA_TEMPR12[49] , \R_DATA_TEMPR12[48] , 
        \R_DATA_TEMPR12[47] , \R_DATA_TEMPR12[46] , 
        \R_DATA_TEMPR12[45] , \R_DATA_TEMPR12[44] , 
        \R_DATA_TEMPR12[43] , \R_DATA_TEMPR12[42] , 
        \R_DATA_TEMPR12[41] , \R_DATA_TEMPR12[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[12][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_1 (.A(\R_DATA_TEMPR8[66] ), .B(\R_DATA_TEMPR9[66] ), .C(
        \R_DATA_TEMPR10[66] ), .D(\R_DATA_TEMPR11[66] ), .Y(OR4_1_Y));
    OR2 OR2_40 (.A(\R_DATA_TEMPR20[20] ), .B(\R_DATA_TEMPR21[20] ), .Y(
        OR2_40_Y));
    OR4 OR4_87 (.A(OR4_151_Y), .B(OR4_554_Y), .C(OR4_98_Y), .D(
        OR4_450_Y), .Y(OR4_87_Y));
    OR4 \OR4_R_DATA[30]  (.A(OR4_37_Y), .B(OR4_214_Y), .C(OR4_529_Y), 
        .D(OR4_264_Y), .Y(R_DATA[30]));
    OR4 OR4_178 (.A(OR4_224_Y), .B(OR4_453_Y), .C(OR4_642_Y), .D(
        OR4_254_Y), .Y(OR4_178_Y));
    OR2 OR2_47 (.A(\R_DATA_TEMPR20[17] ), .B(\R_DATA_TEMPR21[17] ), .Y(
        OR2_47_Y));
    OR4 OR4_159 (.A(\R_DATA_TEMPR8[42] ), .B(\R_DATA_TEMPR9[42] ), .C(
        \R_DATA_TEMPR10[42] ), .D(\R_DATA_TEMPR11[42] ), .Y(OR4_159_Y));
    OR4 OR4_491 (.A(\R_DATA_TEMPR12[11] ), .B(\R_DATA_TEMPR13[11] ), 
        .C(\R_DATA_TEMPR14[11] ), .D(\R_DATA_TEMPR15[11] ), .Y(
        OR4_491_Y));
    OR4 OR4_165 (.A(\R_DATA_TEMPR16[72] ), .B(\R_DATA_TEMPR17[72] ), 
        .C(\R_DATA_TEMPR18[72] ), .D(\R_DATA_TEMPR19[72] ), .Y(
        OR4_165_Y));
    OR4 OR4_133 (.A(OR4_483_Y), .B(OR2_27_Y), .C(\R_DATA_TEMPR22[58] ), 
        .D(\R_DATA_TEMPR23[58] ), .Y(OR4_133_Y));
    OR4 OR4_515 (.A(OR4_140_Y), .B(OR2_19_Y), .C(\R_DATA_TEMPR22[6] ), 
        .D(\R_DATA_TEMPR23[6] ), .Y(OR4_515_Y));
    OR4 OR4_498 (.A(\R_DATA_TEMPR8[73] ), .B(\R_DATA_TEMPR9[73] ), .C(
        \R_DATA_TEMPR10[73] ), .D(\R_DATA_TEMPR11[73] ), .Y(OR4_498_Y));
    OR4 OR4_467 (.A(\R_DATA_TEMPR0[18] ), .B(\R_DATA_TEMPR1[18] ), .C(
        \R_DATA_TEMPR2[18] ), .D(\R_DATA_TEMPR3[18] ), .Y(OR4_467_Y));
    OR4 OR4_92 (.A(\R_DATA_TEMPR0[6] ), .B(\R_DATA_TEMPR1[6] ), .C(
        \R_DATA_TEMPR2[6] ), .D(\R_DATA_TEMPR3[6] ), .Y(OR4_92_Y));
    OR4 \OR4_R_DATA[36]  (.A(OR4_504_Y), .B(OR4_176_Y), .C(OR4_302_Y), 
        .D(OR4_332_Y), .Y(R_DATA[36]));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[1]  (.A(CFG2_6_Y), .B(
        R_ADDR[13]), .C(R_EN), .Y(\BLKY2[1] ));
    OR4 OR4_648 (.A(\R_DATA_TEMPR28[31] ), .B(\R_DATA_TEMPR29[31] ), 
        .C(\R_DATA_TEMPR30[31] ), .D(\R_DATA_TEMPR31[31] ), .Y(
        OR4_648_Y));
    OR4 OR4_685 (.A(\R_DATA_TEMPR0[39] ), .B(\R_DATA_TEMPR1[39] ), .C(
        \R_DATA_TEMPR2[39] ), .D(\R_DATA_TEMPR3[39] ), .Y(OR4_685_Y));
    OR2 OR2_60 (.A(\R_DATA_TEMPR20[64] ), .B(\R_DATA_TEMPR21[64] ), .Y(
        OR2_60_Y));
    OR2 OR2_74 (.A(\R_DATA_TEMPR20[36] ), .B(\R_DATA_TEMPR21[36] ), .Y(
        OR2_74_Y));
    OR4 OR4_613 (.A(\R_DATA_TEMPR12[76] ), .B(\R_DATA_TEMPR13[76] ), 
        .C(\R_DATA_TEMPR14[76] ), .D(\R_DATA_TEMPR15[76] ), .Y(
        OR4_613_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%26%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0 (
        .A_DOUT({\R_DATA_TEMPR26[39] , \R_DATA_TEMPR26[38] , 
        \R_DATA_TEMPR26[37] , \R_DATA_TEMPR26[36] , 
        \R_DATA_TEMPR26[35] , \R_DATA_TEMPR26[34] , 
        \R_DATA_TEMPR26[33] , \R_DATA_TEMPR26[32] , 
        \R_DATA_TEMPR26[31] , \R_DATA_TEMPR26[30] , 
        \R_DATA_TEMPR26[29] , \R_DATA_TEMPR26[28] , 
        \R_DATA_TEMPR26[27] , \R_DATA_TEMPR26[26] , 
        \R_DATA_TEMPR26[25] , \R_DATA_TEMPR26[24] , 
        \R_DATA_TEMPR26[23] , \R_DATA_TEMPR26[22] , 
        \R_DATA_TEMPR26[21] , \R_DATA_TEMPR26[20] }), .B_DOUT({
        \R_DATA_TEMPR26[19] , \R_DATA_TEMPR26[18] , 
        \R_DATA_TEMPR26[17] , \R_DATA_TEMPR26[16] , 
        \R_DATA_TEMPR26[15] , \R_DATA_TEMPR26[14] , 
        \R_DATA_TEMPR26[13] , \R_DATA_TEMPR26[12] , 
        \R_DATA_TEMPR26[11] , \R_DATA_TEMPR26[10] , 
        \R_DATA_TEMPR26[9] , \R_DATA_TEMPR26[8] , \R_DATA_TEMPR26[7] , 
        \R_DATA_TEMPR26[6] , \R_DATA_TEMPR26[5] , \R_DATA_TEMPR26[4] , 
        \R_DATA_TEMPR26[3] , \R_DATA_TEMPR26[2] , \R_DATA_TEMPR26[1] , 
        \R_DATA_TEMPR26[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_642 (.A(\R_DATA_TEMPR8[3] ), .B(\R_DATA_TEMPR9[3] ), .C(
        \R_DATA_TEMPR10[3] ), .D(\R_DATA_TEMPR11[3] ), .Y(OR4_642_Y));
    OR2 OR2_67 (.A(\R_DATA_TEMPR20[16] ), .B(\R_DATA_TEMPR21[16] ), .Y(
        OR2_67_Y));
    CFG2 #( .INIT(4'h8) )  CFG2_0 (.A(W_ADDR[12]), .B(W_ADDR[11]), .Y(
        CFG2_0_Y));
    OR2 OR2_30 (.A(\R_DATA_TEMPR20[35] ), .B(\R_DATA_TEMPR21[35] ), .Y(
        OR2_30_Y));
    OR4 OR4_324 (.A(\R_DATA_TEMPR24[54] ), .B(\R_DATA_TEMPR25[54] ), 
        .C(\R_DATA_TEMPR26[54] ), .D(\R_DATA_TEMPR27[54] ), .Y(
        OR4_324_Y));
    OR4 OR4_265 (.A(OR4_695_Y), .B(OR2_18_Y), .C(\R_DATA_TEMPR22[15] ), 
        .D(\R_DATA_TEMPR23[15] ), .Y(OR4_265_Y));
    OR4 OR4_49 (.A(\R_DATA_TEMPR24[42] ), .B(\R_DATA_TEMPR25[42] ), .C(
        \R_DATA_TEMPR26[42] ), .D(\R_DATA_TEMPR27[42] ), .Y(OR4_49_Y));
    OR4 OR4_599 (.A(OR4_573_Y), .B(OR4_568_Y), .C(OR4_525_Y), .D(
        OR4_702_Y), .Y(OR4_599_Y));
    OR2 OR2_14 (.A(\R_DATA_TEMPR20[32] ), .B(\R_DATA_TEMPR21[32] ), .Y(
        OR2_14_Y));
    OR2 OR2_37 (.A(\R_DATA_TEMPR20[38] ), .B(\R_DATA_TEMPR21[38] ), .Y(
        OR2_37_Y));
    OR4 OR4_590 (.A(\R_DATA_TEMPR4[61] ), .B(\R_DATA_TEMPR5[61] ), .C(
        \R_DATA_TEMPR6[61] ), .D(\R_DATA_TEMPR7[61] ), .Y(OR4_590_Y));
    OR4 OR4_121 (.A(\R_DATA_TEMPR0[36] ), .B(\R_DATA_TEMPR1[36] ), .C(
        \R_DATA_TEMPR2[36] ), .D(\R_DATA_TEMPR3[36] ), .Y(OR4_121_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%30%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0 (
        .A_DOUT({\R_DATA_TEMPR30[39] , \R_DATA_TEMPR30[38] , 
        \R_DATA_TEMPR30[37] , \R_DATA_TEMPR30[36] , 
        \R_DATA_TEMPR30[35] , \R_DATA_TEMPR30[34] , 
        \R_DATA_TEMPR30[33] , \R_DATA_TEMPR30[32] , 
        \R_DATA_TEMPR30[31] , \R_DATA_TEMPR30[30] , 
        \R_DATA_TEMPR30[29] , \R_DATA_TEMPR30[28] , 
        \R_DATA_TEMPR30[27] , \R_DATA_TEMPR30[26] , 
        \R_DATA_TEMPR30[25] , \R_DATA_TEMPR30[24] , 
        \R_DATA_TEMPR30[23] , \R_DATA_TEMPR30[22] , 
        \R_DATA_TEMPR30[21] , \R_DATA_TEMPR30[20] }), .B_DOUT({
        \R_DATA_TEMPR30[19] , \R_DATA_TEMPR30[18] , 
        \R_DATA_TEMPR30[17] , \R_DATA_TEMPR30[16] , 
        \R_DATA_TEMPR30[15] , \R_DATA_TEMPR30[14] , 
        \R_DATA_TEMPR30[13] , \R_DATA_TEMPR30[12] , 
        \R_DATA_TEMPR30[11] , \R_DATA_TEMPR30[10] , 
        \R_DATA_TEMPR30[9] , \R_DATA_TEMPR30[8] , \R_DATA_TEMPR30[7] , 
        \R_DATA_TEMPR30[6] , \R_DATA_TEMPR30[5] , \R_DATA_TEMPR30[4] , 
        \R_DATA_TEMPR30[3] , \R_DATA_TEMPR30[2] , \R_DATA_TEMPR30[1] , 
        \R_DATA_TEMPR30[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR2 OR2_53 (.A(\R_DATA_TEMPR20[65] ), .B(\R_DATA_TEMPR21[65] ), .Y(
        OR2_53_Y));
    OR4 \OR4_R_DATA[18]  (.A(OR4_689_Y), .B(OR4_594_Y), .C(OR4_272_Y), 
        .D(OR4_361_Y), .Y(R_DATA[18]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%3%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C1 (
        .A_DOUT({\R_DATA_TEMPR3[79] , \R_DATA_TEMPR3[78] , 
        \R_DATA_TEMPR3[77] , \R_DATA_TEMPR3[76] , \R_DATA_TEMPR3[75] , 
        \R_DATA_TEMPR3[74] , \R_DATA_TEMPR3[73] , \R_DATA_TEMPR3[72] , 
        \R_DATA_TEMPR3[71] , \R_DATA_TEMPR3[70] , \R_DATA_TEMPR3[69] , 
        \R_DATA_TEMPR3[68] , \R_DATA_TEMPR3[67] , \R_DATA_TEMPR3[66] , 
        \R_DATA_TEMPR3[65] , \R_DATA_TEMPR3[64] , \R_DATA_TEMPR3[63] , 
        \R_DATA_TEMPR3[62] , \R_DATA_TEMPR3[61] , \R_DATA_TEMPR3[60] })
        , .B_DOUT({\R_DATA_TEMPR3[59] , \R_DATA_TEMPR3[58] , 
        \R_DATA_TEMPR3[57] , \R_DATA_TEMPR3[56] , \R_DATA_TEMPR3[55] , 
        \R_DATA_TEMPR3[54] , \R_DATA_TEMPR3[53] , \R_DATA_TEMPR3[52] , 
        \R_DATA_TEMPR3[51] , \R_DATA_TEMPR3[50] , \R_DATA_TEMPR3[49] , 
        \R_DATA_TEMPR3[48] , \R_DATA_TEMPR3[47] , \R_DATA_TEMPR3[46] , 
        \R_DATA_TEMPR3[45] , \R_DATA_TEMPR3[44] , \R_DATA_TEMPR3[43] , 
        \R_DATA_TEMPR3[42] , \R_DATA_TEMPR3[41] , \R_DATA_TEMPR3[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[3][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[0] , 
        R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[0] , W_ADDR[10], W_ADDR[9]}), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_680 (.A(OR4_99_Y), .B(OR2_69_Y), .C(\R_DATA_TEMPR22[0] ), 
        .D(\R_DATA_TEMPR23[0] ), .Y(OR4_680_Y));
    OR4 OR4_113 (.A(\R_DATA_TEMPR16[13] ), .B(\R_DATA_TEMPR17[13] ), 
        .C(\R_DATA_TEMPR18[13] ), .D(\R_DATA_TEMPR19[13] ), .Y(
        OR4_113_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%1%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C1 (
        .A_DOUT({\R_DATA_TEMPR1[79] , \R_DATA_TEMPR1[78] , 
        \R_DATA_TEMPR1[77] , \R_DATA_TEMPR1[76] , \R_DATA_TEMPR1[75] , 
        \R_DATA_TEMPR1[74] , \R_DATA_TEMPR1[73] , \R_DATA_TEMPR1[72] , 
        \R_DATA_TEMPR1[71] , \R_DATA_TEMPR1[70] , \R_DATA_TEMPR1[69] , 
        \R_DATA_TEMPR1[68] , \R_DATA_TEMPR1[67] , \R_DATA_TEMPR1[66] , 
        \R_DATA_TEMPR1[65] , \R_DATA_TEMPR1[64] , \R_DATA_TEMPR1[63] , 
        \R_DATA_TEMPR1[62] , \R_DATA_TEMPR1[61] , \R_DATA_TEMPR1[60] })
        , .B_DOUT({\R_DATA_TEMPR1[59] , \R_DATA_TEMPR1[58] , 
        \R_DATA_TEMPR1[57] , \R_DATA_TEMPR1[56] , \R_DATA_TEMPR1[55] , 
        \R_DATA_TEMPR1[54] , \R_DATA_TEMPR1[53] , \R_DATA_TEMPR1[52] , 
        \R_DATA_TEMPR1[51] , \R_DATA_TEMPR1[50] , \R_DATA_TEMPR1[49] , 
        \R_DATA_TEMPR1[48] , \R_DATA_TEMPR1[47] , \R_DATA_TEMPR1[46] , 
        \R_DATA_TEMPR1[45] , \R_DATA_TEMPR1[44] , \R_DATA_TEMPR1[43] , 
        \R_DATA_TEMPR1[42] , \R_DATA_TEMPR1[41] , \R_DATA_TEMPR1[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[1][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[0] , 
        \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_132 (.A(\R_DATA_TEMPR8[28] ), .B(\R_DATA_TEMPR9[28] ), .C(
        \R_DATA_TEMPR10[28] ), .D(\R_DATA_TEMPR11[28] ), .Y(OR4_132_Y));
    OR4 OR4_7 (.A(\R_DATA_TEMPR4[79] ), .B(\R_DATA_TEMPR5[79] ), .C(
        \R_DATA_TEMPR6[79] ), .D(\R_DATA_TEMPR7[79] ), .Y(OR4_7_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%11%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C1 (
        .A_DOUT({\R_DATA_TEMPR11[79] , \R_DATA_TEMPR11[78] , 
        \R_DATA_TEMPR11[77] , \R_DATA_TEMPR11[76] , 
        \R_DATA_TEMPR11[75] , \R_DATA_TEMPR11[74] , 
        \R_DATA_TEMPR11[73] , \R_DATA_TEMPR11[72] , 
        \R_DATA_TEMPR11[71] , \R_DATA_TEMPR11[70] , 
        \R_DATA_TEMPR11[69] , \R_DATA_TEMPR11[68] , 
        \R_DATA_TEMPR11[67] , \R_DATA_TEMPR11[66] , 
        \R_DATA_TEMPR11[65] , \R_DATA_TEMPR11[64] , 
        \R_DATA_TEMPR11[63] , \R_DATA_TEMPR11[62] , 
        \R_DATA_TEMPR11[61] , \R_DATA_TEMPR11[60] }), .B_DOUT({
        \R_DATA_TEMPR11[59] , \R_DATA_TEMPR11[58] , 
        \R_DATA_TEMPR11[57] , \R_DATA_TEMPR11[56] , 
        \R_DATA_TEMPR11[55] , \R_DATA_TEMPR11[54] , 
        \R_DATA_TEMPR11[53] , \R_DATA_TEMPR11[52] , 
        \R_DATA_TEMPR11[51] , \R_DATA_TEMPR11[50] , 
        \R_DATA_TEMPR11[49] , \R_DATA_TEMPR11[48] , 
        \R_DATA_TEMPR11[47] , \R_DATA_TEMPR11[46] , 
        \R_DATA_TEMPR11[45] , \R_DATA_TEMPR11[44] , 
        \R_DATA_TEMPR11[43] , \R_DATA_TEMPR11[42] , 
        \R_DATA_TEMPR11[41] , \R_DATA_TEMPR11[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[11][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_421 (.A(OR4_484_Y), .B(OR4_158_Y), .C(OR4_429_Y), .D(
        OR4_55_Y), .Y(OR4_421_Y));
    OR4 OR4_463 (.A(\R_DATA_TEMPR12[4] ), .B(\R_DATA_TEMPR13[4] ), .C(
        \R_DATA_TEMPR14[4] ), .D(\R_DATA_TEMPR15[4] ), .Y(OR4_463_Y));
    OR4 OR4_661 (.A(OR4_211_Y), .B(OR2_49_Y), .C(\R_DATA_TEMPR22[7] ), 
        .D(\R_DATA_TEMPR23[7] ), .Y(OR4_661_Y));
    OR4 OR4_657 (.A(\R_DATA_TEMPR24[77] ), .B(\R_DATA_TEMPR25[77] ), 
        .C(\R_DATA_TEMPR26[77] ), .D(\R_DATA_TEMPR27[77] ), .Y(
        OR4_657_Y));
    OR4 OR4_428 (.A(OR4_631_Y), .B(OR2_28_Y), .C(\R_DATA_TEMPR22[14] ), 
        .D(\R_DATA_TEMPR23[14] ), .Y(OR4_428_Y));
    OR4 OR4_268 (.A(\R_DATA_TEMPR4[28] ), .B(\R_DATA_TEMPR5[28] ), .C(
        \R_DATA_TEMPR6[28] ), .D(\R_DATA_TEMPR7[28] ), .Y(OR4_268_Y));
    OR4 OR4_387 (.A(\R_DATA_TEMPR8[8] ), .B(\R_DATA_TEMPR9[8] ), .C(
        \R_DATA_TEMPR10[8] ), .D(\R_DATA_TEMPR11[8] ), .Y(OR4_387_Y));
    OR4 OR4_180 (.A(\R_DATA_TEMPR28[73] ), .B(\R_DATA_TEMPR29[73] ), 
        .C(\R_DATA_TEMPR30[73] ), .D(\R_DATA_TEMPR31[73] ), .Y(
        OR4_180_Y));
    OR4 OR4_105 (.A(\R_DATA_TEMPR16[5] ), .B(\R_DATA_TEMPR17[5] ), .C(
        \R_DATA_TEMPR18[5] ), .D(\R_DATA_TEMPR19[5] ), .Y(OR4_105_Y));
    OR4 OR4_407 (.A(\R_DATA_TEMPR4[26] ), .B(\R_DATA_TEMPR5[26] ), .C(
        \R_DATA_TEMPR6[26] ), .D(\R_DATA_TEMPR7[26] ), .Y(OR4_407_Y));
    OR4 OR4_175 (.A(\R_DATA_TEMPR16[54] ), .B(\R_DATA_TEMPR17[54] ), 
        .C(\R_DATA_TEMPR18[54] ), .D(\R_DATA_TEMPR19[54] ), .Y(
        OR4_175_Y));
    OR4 OR4_393 (.A(OR4_685_Y), .B(OR4_221_Y), .C(OR4_519_Y), .D(
        OR4_85_Y), .Y(OR4_393_Y));
    OR4 OR4_239 (.A(\R_DATA_TEMPR0[9] ), .B(\R_DATA_TEMPR1[9] ), .C(
        \R_DATA_TEMPR2[9] ), .D(\R_DATA_TEMPR3[9] ), .Y(OR4_239_Y));
    OR4 OR4_42 (.A(OR4_357_Y), .B(OR2_33_Y), .C(\R_DATA_TEMPR22[79] ), 
        .D(\R_DATA_TEMPR23[79] ), .Y(OR4_42_Y));
    OR4 OR4_529 (.A(\R_DATA_TEMPR24[30] ), .B(\R_DATA_TEMPR25[30] ), 
        .C(\R_DATA_TEMPR26[30] ), .D(\R_DATA_TEMPR27[30] ), .Y(
        OR4_529_Y));
    OR4 OR4_477 (.A(\R_DATA_TEMPR4[23] ), .B(\R_DATA_TEMPR5[23] ), .C(
        \R_DATA_TEMPR6[23] ), .D(\R_DATA_TEMPR7[23] ), .Y(OR4_477_Y));
    OR4 OR4_492 (.A(\R_DATA_TEMPR0[79] ), .B(\R_DATA_TEMPR1[79] ), .C(
        \R_DATA_TEMPR2[79] ), .D(\R_DATA_TEMPR3[79] ), .Y(OR4_492_Y));
    OR4 OR4_520 (.A(OR4_251_Y), .B(OR2_17_Y), .C(\R_DATA_TEMPR22[55] ), 
        .D(\R_DATA_TEMPR23[55] ), .Y(OR4_520_Y));
    OR2 OR2_51 (.A(\R_DATA_TEMPR20[24] ), .B(\R_DATA_TEMPR21[24] ), .Y(
        OR2_51_Y));
    OR4 OR4_499 (.A(\R_DATA_TEMPR24[2] ), .B(\R_DATA_TEMPR25[2] ), .C(
        \R_DATA_TEMPR26[2] ), .D(\R_DATA_TEMPR27[2] ), .Y(OR4_499_Y));
    OR4 OR4_88 (.A(OR4_325_Y), .B(OR4_201_Y), .C(OR4_185_Y), .D(
        OR4_620_Y), .Y(OR4_88_Y));
    OR4 OR4_205 (.A(OR4_637_Y), .B(OR2_44_Y), .C(\R_DATA_TEMPR22[25] ), 
        .D(\R_DATA_TEMPR23[25] ), .Y(OR4_205_Y));
    OR4 OR4_188 (.A(\R_DATA_TEMPR0[66] ), .B(\R_DATA_TEMPR1[66] ), .C(
        \R_DATA_TEMPR2[66] ), .D(\R_DATA_TEMPR3[66] ), .Y(OR4_188_Y));
    OR4 OR4_196 (.A(\R_DATA_TEMPR8[55] ), .B(\R_DATA_TEMPR9[55] ), .C(
        \R_DATA_TEMPR10[55] ), .D(\R_DATA_TEMPR11[55] ), .Y(OR4_196_Y));
    OR4 OR4_112 (.A(\R_DATA_TEMPR16[64] ), .B(\R_DATA_TEMPR17[64] ), 
        .C(\R_DATA_TEMPR18[64] ), .D(\R_DATA_TEMPR19[64] ), .Y(
        OR4_112_Y));
    OR2 OR2_48 (.A(\R_DATA_TEMPR20[49] ), .B(\R_DATA_TEMPR21[49] ), .Y(
        OR2_48_Y));
    OR4 \OR4_R_DATA[48]  (.A(OR4_338_Y), .B(OR4_258_Y), .C(OR4_641_Y), 
        .D(OR4_13_Y), .Y(R_DATA[48]));
    OR4 OR4_275 (.A(\R_DATA_TEMPR24[8] ), .B(\R_DATA_TEMPR25[8] ), .C(
        \R_DATA_TEMPR26[8] ), .D(\R_DATA_TEMPR27[8] ), .Y(OR4_275_Y));
    OR4 OR4_646 (.A(\R_DATA_TEMPR8[15] ), .B(\R_DATA_TEMPR9[15] ), .C(
        \R_DATA_TEMPR10[15] ), .D(\R_DATA_TEMPR11[15] ), .Y(OR4_646_Y));
    OR4 \OR4_R_DATA[37]  (.A(OR4_316_Y), .B(OR4_670_Y), .C(OR4_119_Y), 
        .D(OR4_208_Y), .Y(R_DATA[37]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%25%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C1 (
        .A_DOUT({\R_DATA_TEMPR25[79] , \R_DATA_TEMPR25[78] , 
        \R_DATA_TEMPR25[77] , \R_DATA_TEMPR25[76] , 
        \R_DATA_TEMPR25[75] , \R_DATA_TEMPR25[74] , 
        \R_DATA_TEMPR25[73] , \R_DATA_TEMPR25[72] , 
        \R_DATA_TEMPR25[71] , \R_DATA_TEMPR25[70] , 
        \R_DATA_TEMPR25[69] , \R_DATA_TEMPR25[68] , 
        \R_DATA_TEMPR25[67] , \R_DATA_TEMPR25[66] , 
        \R_DATA_TEMPR25[65] , \R_DATA_TEMPR25[64] , 
        \R_DATA_TEMPR25[63] , \R_DATA_TEMPR25[62] , 
        \R_DATA_TEMPR25[61] , \R_DATA_TEMPR25[60] }), .B_DOUT({
        \R_DATA_TEMPR25[59] , \R_DATA_TEMPR25[58] , 
        \R_DATA_TEMPR25[57] , \R_DATA_TEMPR25[56] , 
        \R_DATA_TEMPR25[55] , \R_DATA_TEMPR25[54] , 
        \R_DATA_TEMPR25[53] , \R_DATA_TEMPR25[52] , 
        \R_DATA_TEMPR25[51] , \R_DATA_TEMPR25[50] , 
        \R_DATA_TEMPR25[49] , \R_DATA_TEMPR25[48] , 
        \R_DATA_TEMPR25[47] , \R_DATA_TEMPR25[46] , 
        \R_DATA_TEMPR25[45] , \R_DATA_TEMPR25[44] , 
        \R_DATA_TEMPR25[43] , \R_DATA_TEMPR25[42] , 
        \R_DATA_TEMPR25[41] , \R_DATA_TEMPR25[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[25][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_257 (.A(\R_DATA_TEMPR28[67] ), .B(\R_DATA_TEMPR29[67] ), 
        .C(\R_DATA_TEMPR30[67] ), .D(\R_DATA_TEMPR31[67] ), .Y(
        OR4_257_Y));
    OR4 OR4_398 (.A(\R_DATA_TEMPR24[12] ), .B(\R_DATA_TEMPR25[12] ), 
        .C(\R_DATA_TEMPR26[12] ), .D(\R_DATA_TEMPR27[12] ), .Y(
        OR4_398_Y));
    OR4 OR4_157 (.A(\R_DATA_TEMPR12[9] ), .B(\R_DATA_TEMPR13[9] ), .C(
        \R_DATA_TEMPR14[9] ), .D(\R_DATA_TEMPR15[9] ), .Y(OR4_157_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%5%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C1 (
        .A_DOUT({\R_DATA_TEMPR5[79] , \R_DATA_TEMPR5[78] , 
        \R_DATA_TEMPR5[77] , \R_DATA_TEMPR5[76] , \R_DATA_TEMPR5[75] , 
        \R_DATA_TEMPR5[74] , \R_DATA_TEMPR5[73] , \R_DATA_TEMPR5[72] , 
        \R_DATA_TEMPR5[71] , \R_DATA_TEMPR5[70] , \R_DATA_TEMPR5[69] , 
        \R_DATA_TEMPR5[68] , \R_DATA_TEMPR5[67] , \R_DATA_TEMPR5[66] , 
        \R_DATA_TEMPR5[65] , \R_DATA_TEMPR5[64] , \R_DATA_TEMPR5[63] , 
        \R_DATA_TEMPR5[62] , \R_DATA_TEMPR5[61] , \R_DATA_TEMPR5[60] })
        , .B_DOUT({\R_DATA_TEMPR5[59] , \R_DATA_TEMPR5[58] , 
        \R_DATA_TEMPR5[57] , \R_DATA_TEMPR5[56] , \R_DATA_TEMPR5[55] , 
        \R_DATA_TEMPR5[54] , \R_DATA_TEMPR5[53] , \R_DATA_TEMPR5[52] , 
        \R_DATA_TEMPR5[51] , \R_DATA_TEMPR5[50] , \R_DATA_TEMPR5[49] , 
        \R_DATA_TEMPR5[48] , \R_DATA_TEMPR5[47] , \R_DATA_TEMPR5[46] , 
        \R_DATA_TEMPR5[45] , \R_DATA_TEMPR5[44] , \R_DATA_TEMPR5[43] , 
        \R_DATA_TEMPR5[42] , \R_DATA_TEMPR5[41] , \R_DATA_TEMPR5[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[5][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[1] , 
        \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_561 (.A(\R_DATA_TEMPR28[29] ), .B(\R_DATA_TEMPR29[29] ), 
        .C(\R_DATA_TEMPR30[29] ), .D(\R_DATA_TEMPR31[29] ), .Y(
        OR4_561_Y));
    OR4 OR4_403 (.A(OR4_518_Y), .B(OR2_5_Y), .C(\R_DATA_TEMPR22[40] ), 
        .D(\R_DATA_TEMPR23[40] ), .Y(OR4_403_Y));
    OR4 OR4_601 (.A(\R_DATA_TEMPR28[5] ), .B(\R_DATA_TEMPR29[5] ), .C(
        \R_DATA_TEMPR30[5] ), .D(\R_DATA_TEMPR31[5] ), .Y(OR4_601_Y));
    OR2 OR2_68 (.A(\R_DATA_TEMPR20[1] ), .B(\R_DATA_TEMPR21[1] ), .Y(
        OR2_68_Y));
    OR4 OR4_208 (.A(\R_DATA_TEMPR28[37] ), .B(\R_DATA_TEMPR29[37] ), 
        .C(\R_DATA_TEMPR30[37] ), .D(\R_DATA_TEMPR31[37] ), .Y(
        OR4_208_Y));
    OR4 OR4_219 (.A(\R_DATA_TEMPR28[13] ), .B(\R_DATA_TEMPR29[13] ), 
        .C(\R_DATA_TEMPR30[13] ), .D(\R_DATA_TEMPR31[13] ), .Y(
        OR4_219_Y));
    OR4 OR4_323 (.A(\R_DATA_TEMPR24[70] ), .B(\R_DATA_TEMPR25[70] ), 
        .C(\R_DATA_TEMPR26[70] ), .D(\R_DATA_TEMPR27[70] ), .Y(
        OR4_323_Y));
    OR4 \OR4_R_DATA[68]  (.A(OR4_191_Y), .B(OR4_83_Y), .C(OR4_482_Y), 
        .D(OR4_580_Y), .Y(R_DATA[68]));
    OR4 \OR4_R_DATA[19]  (.A(OR4_240_Y), .B(OR4_66_Y), .C(OR4_24_Y), 
        .D(OR4_621_Y), .Y(R_DATA[19]));
    OR4 OR4_473 (.A(OR4_370_Y), .B(OR2_23_Y), .C(\R_DATA_TEMPR22[77] ), 
        .D(\R_DATA_TEMPR23[77] ), .Y(OR4_473_Y));
    OR4 OR4_671 (.A(\R_DATA_TEMPR24[52] ), .B(\R_DATA_TEMPR25[52] ), 
        .C(\R_DATA_TEMPR26[52] ), .D(\R_DATA_TEMPR27[52] ), .Y(
        OR4_671_Y));
    OR2 OR2_38 (.A(\R_DATA_TEMPR20[47] ), .B(\R_DATA_TEMPR21[47] ), .Y(
        OR2_38_Y));
    OR4 \OR4_R_DATA[75]  (.A(OR4_605_Y), .B(OR4_234_Y), .C(OR4_505_Y), 
        .D(OR4_298_Y), .Y(R_DATA[75]));
    OR4 OR4_422 (.A(OR4_696_Y), .B(OR4_96_Y), .C(OR4_533_Y), .D(
        OR4_443_Y), .Y(OR4_422_Y));
    OR4 OR4_278 (.A(\R_DATA_TEMPR28[49] ), .B(\R_DATA_TEMPR29[49] ), 
        .C(\R_DATA_TEMPR30[49] ), .D(\R_DATA_TEMPR31[49] ), .Y(
        OR4_278_Y));
    OR4 OR4_23 (.A(\R_DATA_TEMPR4[41] ), .B(\R_DATA_TEMPR5[41] ), .C(
        \R_DATA_TEMPR6[41] ), .D(\R_DATA_TEMPR7[41] ), .Y(OR4_23_Y));
    OR4 OR4_199 (.A(\R_DATA_TEMPR0[40] ), .B(\R_DATA_TEMPR1[40] ), .C(
        \R_DATA_TEMPR2[40] ), .D(\R_DATA_TEMPR3[40] ), .Y(OR4_199_Y));
    OR4 OR4_254 (.A(\R_DATA_TEMPR12[3] ), .B(\R_DATA_TEMPR13[3] ), .C(
        \R_DATA_TEMPR14[3] ), .D(\R_DATA_TEMPR15[3] ), .Y(OR4_254_Y));
    OR4 OR4_429 (.A(\R_DATA_TEMPR8[57] ), .B(\R_DATA_TEMPR9[57] ), .C(
        \R_DATA_TEMPR10[57] ), .D(\R_DATA_TEMPR11[57] ), .Y(OR4_429_Y));
    OR4 OR4_262 (.A(\R_DATA_TEMPR0[11] ), .B(\R_DATA_TEMPR1[11] ), .C(
        \R_DATA_TEMPR2[11] ), .D(\R_DATA_TEMPR3[11] ), .Y(OR4_262_Y));
    OR4 OR4_126 (.A(OR4_345_Y), .B(OR2_39_Y), .C(\R_DATA_TEMPR22[31] ), 
        .D(\R_DATA_TEMPR23[31] ), .Y(OR4_126_Y));
    OR4 OR4_94 (.A(\R_DATA_TEMPR4[65] ), .B(\R_DATA_TEMPR5[65] ), .C(
        \R_DATA_TEMPR6[65] ), .D(\R_DATA_TEMPR7[65] ), .Y(OR4_94_Y));
    OR4 OR4_65 (.A(\R_DATA_TEMPR16[34] ), .B(\R_DATA_TEMPR17[34] ), .C(
        \R_DATA_TEMPR18[34] ), .D(\R_DATA_TEMPR19[34] ), .Y(OR4_65_Y));
    OR4 OR4_360 (.A(\R_DATA_TEMPR16[32] ), .B(\R_DATA_TEMPR17[32] ), 
        .C(\R_DATA_TEMPR18[32] ), .D(\R_DATA_TEMPR19[32] ), .Y(
        OR4_360_Y));
    OR4 OR4_355 (.A(\R_DATA_TEMPR16[60] ), .B(\R_DATA_TEMPR17[60] ), 
        .C(\R_DATA_TEMPR18[60] ), .D(\R_DATA_TEMPR19[60] ), .Y(
        OR4_355_Y));
    OR4 OR4_328 (.A(\R_DATA_TEMPR8[37] ), .B(\R_DATA_TEMPR9[37] ), .C(
        \R_DATA_TEMPR10[37] ), .D(\R_DATA_TEMPR11[37] ), .Y(OR4_328_Y));
    OR4 OR4_344 (.A(\R_DATA_TEMPR28[52] ), .B(\R_DATA_TEMPR29[52] ), 
        .C(\R_DATA_TEMPR30[52] ), .D(\R_DATA_TEMPR31[52] ), .Y(
        OR4_344_Y));
    OR4 OR4_185 (.A(\R_DATA_TEMPR8[43] ), .B(\R_DATA_TEMPR9[43] ), .C(
        \R_DATA_TEMPR10[43] ), .D(\R_DATA_TEMPR11[43] ), .Y(OR4_185_Y));
    OR4 OR4_141 (.A(\R_DATA_TEMPR28[76] ), .B(\R_DATA_TEMPR29[76] ), 
        .C(\R_DATA_TEMPR30[76] ), .D(\R_DATA_TEMPR31[76] ), .Y(
        OR4_141_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%25%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0 (
        .A_DOUT({\R_DATA_TEMPR25[39] , \R_DATA_TEMPR25[38] , 
        \R_DATA_TEMPR25[37] , \R_DATA_TEMPR25[36] , 
        \R_DATA_TEMPR25[35] , \R_DATA_TEMPR25[34] , 
        \R_DATA_TEMPR25[33] , \R_DATA_TEMPR25[32] , 
        \R_DATA_TEMPR25[31] , \R_DATA_TEMPR25[30] , 
        \R_DATA_TEMPR25[29] , \R_DATA_TEMPR25[28] , 
        \R_DATA_TEMPR25[27] , \R_DATA_TEMPR25[26] , 
        \R_DATA_TEMPR25[25] , \R_DATA_TEMPR25[24] , 
        \R_DATA_TEMPR25[23] , \R_DATA_TEMPR25[22] , 
        \R_DATA_TEMPR25[21] , \R_DATA_TEMPR25[20] }), .B_DOUT({
        \R_DATA_TEMPR25[19] , \R_DATA_TEMPR25[18] , 
        \R_DATA_TEMPR25[17] , \R_DATA_TEMPR25[16] , 
        \R_DATA_TEMPR25[15] , \R_DATA_TEMPR25[14] , 
        \R_DATA_TEMPR25[13] , \R_DATA_TEMPR25[12] , 
        \R_DATA_TEMPR25[11] , \R_DATA_TEMPR25[10] , 
        \R_DATA_TEMPR25[9] , \R_DATA_TEMPR25[8] , \R_DATA_TEMPR25[7] , 
        \R_DATA_TEMPR25[6] , \R_DATA_TEMPR25[5] , \R_DATA_TEMPR25[4] , 
        \R_DATA_TEMPR25[3] , \R_DATA_TEMPR25[2] , \R_DATA_TEMPR25[1] , 
        \R_DATA_TEMPR25[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_717 (.A(\R_DATA_TEMPR28[77] ), .B(\R_DATA_TEMPR29[77] ), 
        .C(\R_DATA_TEMPR30[77] ), .D(\R_DATA_TEMPR31[77] ), .Y(
        OR4_717_Y));
    OR4 \OR4_R_DATA[49]  (.A(OR4_607_Y), .B(OR4_440_Y), .C(OR4_395_Y), 
        .D(OR4_278_Y), .Y(R_DATA[49]));
    OR4 OR4_36 (.A(\R_DATA_TEMPR8[60] ), .B(\R_DATA_TEMPR9[60] ), .C(
        \R_DATA_TEMPR10[60] ), .D(\R_DATA_TEMPR11[60] ), .Y(OR4_36_Y));
    OR4 OR4_487 (.A(\R_DATA_TEMPR8[76] ), .B(\R_DATA_TEMPR9[76] ), .C(
        \R_DATA_TEMPR10[76] ), .D(\R_DATA_TEMPR11[76] ), .Y(OR4_487_Y));
    OR4 OR4_714 (.A(\R_DATA_TEMPR24[79] ), .B(\R_DATA_TEMPR25[79] ), 
        .C(\R_DATA_TEMPR26[79] ), .D(\R_DATA_TEMPR27[79] ), .Y(
        OR4_714_Y));
    OR4 OR4_501 (.A(OR4_397_Y), .B(OR2_47_Y), .C(\R_DATA_TEMPR22[17] ), 
        .D(\R_DATA_TEMPR23[17] ), .Y(OR4_501_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%27%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0 (
        .A_DOUT({\R_DATA_TEMPR27[39] , \R_DATA_TEMPR27[38] , 
        \R_DATA_TEMPR27[37] , \R_DATA_TEMPR27[36] , 
        \R_DATA_TEMPR27[35] , \R_DATA_TEMPR27[34] , 
        \R_DATA_TEMPR27[33] , \R_DATA_TEMPR27[32] , 
        \R_DATA_TEMPR27[31] , \R_DATA_TEMPR27[30] , 
        \R_DATA_TEMPR27[29] , \R_DATA_TEMPR27[28] , 
        \R_DATA_TEMPR27[27] , \R_DATA_TEMPR27[26] , 
        \R_DATA_TEMPR27[25] , \R_DATA_TEMPR27[24] , 
        \R_DATA_TEMPR27[23] , \R_DATA_TEMPR27[22] , 
        \R_DATA_TEMPR27[21] , \R_DATA_TEMPR27[20] }), .B_DOUT({
        \R_DATA_TEMPR27[19] , \R_DATA_TEMPR27[18] , 
        \R_DATA_TEMPR27[17] , \R_DATA_TEMPR27[16] , 
        \R_DATA_TEMPR27[15] , \R_DATA_TEMPR27[14] , 
        \R_DATA_TEMPR27[13] , \R_DATA_TEMPR27[12] , 
        \R_DATA_TEMPR27[11] , \R_DATA_TEMPR27[10] , 
        \R_DATA_TEMPR27[9] , \R_DATA_TEMPR27[8] , \R_DATA_TEMPR27[7] , 
        \R_DATA_TEMPR27[6] , \R_DATA_TEMPR27[5] , \R_DATA_TEMPR27[4] , 
        \R_DATA_TEMPR27[3] , \R_DATA_TEMPR27[2] , \R_DATA_TEMPR27[1] , 
        \R_DATA_TEMPR27[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_21 (.A(\R_DATA_TEMPR8[63] ), .B(\R_DATA_TEMPR9[63] ), .C(
        \R_DATA_TEMPR10[63] ), .D(\R_DATA_TEMPR11[63] ), .Y(OR4_21_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[3]  (.A(CFG2_5_Y), .B(
        R_ADDR[13]), .C(R_EN), .Y(\BLKY2[3] ));
    OR4 OR4_129 (.A(\R_DATA_TEMPR24[16] ), .B(\R_DATA_TEMPR25[16] ), 
        .C(\R_DATA_TEMPR26[16] ), .D(\R_DATA_TEMPR27[16] ), .Y(
        OR4_129_Y));
    OR4 OR4_571 (.A(OR4_123_Y), .B(OR4_552_Y), .C(OR4_582_Y), .D(
        OR4_237_Y), .Y(OR4_571_Y));
    OR4 OR4_441 (.A(OR4_479_Y), .B(OR2_42_Y), .C(\R_DATA_TEMPR22[8] ), 
        .D(\R_DATA_TEMPR23[8] ), .Y(OR4_441_Y));
    OR4 OR4_697 (.A(\R_DATA_TEMPR28[61] ), .B(\R_DATA_TEMPR29[61] ), 
        .C(\R_DATA_TEMPR30[61] ), .D(\R_DATA_TEMPR31[61] ), .Y(
        OR4_697_Y));
    OR4 OR4_448 (.A(\R_DATA_TEMPR28[42] ), .B(\R_DATA_TEMPR29[42] ), 
        .C(\R_DATA_TEMPR30[42] ), .D(\R_DATA_TEMPR31[42] ), .Y(
        OR4_448_Y));
    OR4 OR4_285 (.A(\R_DATA_TEMPR16[33] ), .B(\R_DATA_TEMPR17[33] ), 
        .C(\R_DATA_TEMPR18[33] ), .D(\R_DATA_TEMPR19[33] ), .Y(
        OR4_285_Y));
    OR4 OR4_202 (.A(\R_DATA_TEMPR24[39] ), .B(\R_DATA_TEMPR25[39] ), 
        .C(\R_DATA_TEMPR26[39] ), .D(\R_DATA_TEMPR27[39] ), .Y(
        OR4_202_Y));
    OR4 OR4_655 (.A(\R_DATA_TEMPR16[59] ), .B(\R_DATA_TEMPR17[59] ), 
        .C(\R_DATA_TEMPR18[59] ), .D(\R_DATA_TEMPR19[59] ), .Y(
        OR4_655_Y));
    OR4 \OR4_R_DATA[69]  (.A(OR4_439_Y), .B(OR4_286_Y), .C(OR4_253_Y), 
        .D(OR4_103_Y), .Y(R_DATA[69]));
    OR4 OR4_272 (.A(\R_DATA_TEMPR24[18] ), .B(\R_DATA_TEMPR25[18] ), 
        .C(\R_DATA_TEMPR26[18] ), .D(\R_DATA_TEMPR27[18] ), .Y(
        OR4_272_Y));
    OR4 OR4_565 (.A(\R_DATA_TEMPR0[45] ), .B(\R_DATA_TEMPR1[45] ), .C(
        \R_DATA_TEMPR2[45] ), .D(\R_DATA_TEMPR3[45] ), .Y(OR4_565_Y));
    OR4 OR4_44 (.A(OR4_461_Y), .B(OR2_2_Y), .C(\R_DATA_TEMPR22[52] ), 
        .D(\R_DATA_TEMPR23[52] ), .Y(OR4_44_Y));
    OR4 OR4_549 (.A(\R_DATA_TEMPR4[30] ), .B(\R_DATA_TEMPR5[30] ), .C(
        \R_DATA_TEMPR6[30] ), .D(\R_DATA_TEMPR7[30] ), .Y(OR4_549_Y));
    OR4 OR4_435 (.A(\R_DATA_TEMPR24[63] ), .B(\R_DATA_TEMPR25[63] ), 
        .C(\R_DATA_TEMPR26[63] ), .D(\R_DATA_TEMPR27[63] ), .Y(
        OR4_435_Y));
    OR4 OR4_300 (.A(OR4_406_Y), .B(OR2_11_Y), .C(\R_DATA_TEMPR22[50] ), 
        .D(\R_DATA_TEMPR23[50] ), .Y(OR4_300_Y));
    OR4 OR4_540 (.A(\R_DATA_TEMPR4[31] ), .B(\R_DATA_TEMPR5[31] ), .C(
        \R_DATA_TEMPR6[31] ), .D(\R_DATA_TEMPR7[31] ), .Y(OR4_540_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[0]  (.A(CFG2_4_Y), .B(
        W_ADDR[13]), .C(W_EN), .Y(\BLKX2[0] ));
    OR4 OR4_483 (.A(\R_DATA_TEMPR16[58] ), .B(\R_DATA_TEMPR17[58] ), 
        .C(\R_DATA_TEMPR18[58] ), .D(\R_DATA_TEMPR19[58] ), .Y(
        OR4_483_Y));
    OR4 OR4_681 (.A(\R_DATA_TEMPR24[29] ), .B(\R_DATA_TEMPR25[29] ), 
        .C(\R_DATA_TEMPR26[29] ), .D(\R_DATA_TEMPR27[29] ), .Y(
        OR4_681_Y));
    OR4 OR4_663 (.A(\R_DATA_TEMPR12[45] ), .B(\R_DATA_TEMPR13[45] ), 
        .C(\R_DATA_TEMPR14[45] ), .D(\R_DATA_TEMPR15[45] ), .Y(
        OR4_663_Y));
    OR4 OR4_370 (.A(\R_DATA_TEMPR16[77] ), .B(\R_DATA_TEMPR17[77] ), 
        .C(\R_DATA_TEMPR18[77] ), .D(\R_DATA_TEMPR19[77] ), .Y(
        OR4_370_Y));
    OR4 OR4_288 (.A(\R_DATA_TEMPR8[29] ), .B(\R_DATA_TEMPR9[29] ), .C(
        \R_DATA_TEMPR10[29] ), .D(\R_DATA_TEMPR11[29] ), .Y(OR4_288_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%29%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C1 (
        .A_DOUT({\R_DATA_TEMPR29[79] , \R_DATA_TEMPR29[78] , 
        \R_DATA_TEMPR29[77] , \R_DATA_TEMPR29[76] , 
        \R_DATA_TEMPR29[75] , \R_DATA_TEMPR29[74] , 
        \R_DATA_TEMPR29[73] , \R_DATA_TEMPR29[72] , 
        \R_DATA_TEMPR29[71] , \R_DATA_TEMPR29[70] , 
        \R_DATA_TEMPR29[69] , \R_DATA_TEMPR29[68] , 
        \R_DATA_TEMPR29[67] , \R_DATA_TEMPR29[66] , 
        \R_DATA_TEMPR29[65] , \R_DATA_TEMPR29[64] , 
        \R_DATA_TEMPR29[63] , \R_DATA_TEMPR29[62] , 
        \R_DATA_TEMPR29[61] , \R_DATA_TEMPR29[60] }), .B_DOUT({
        \R_DATA_TEMPR29[59] , \R_DATA_TEMPR29[58] , 
        \R_DATA_TEMPR29[57] , \R_DATA_TEMPR29[56] , 
        \R_DATA_TEMPR29[55] , \R_DATA_TEMPR29[54] , 
        \R_DATA_TEMPR29[53] , \R_DATA_TEMPR29[52] , 
        \R_DATA_TEMPR29[51] , \R_DATA_TEMPR29[50] , 
        \R_DATA_TEMPR29[49] , \R_DATA_TEMPR29[48] , 
        \R_DATA_TEMPR29[47] , \R_DATA_TEMPR29[46] , 
        \R_DATA_TEMPR29[45] , \R_DATA_TEMPR29[44] , 
        \R_DATA_TEMPR29[43] , \R_DATA_TEMPR29[42] , 
        \R_DATA_TEMPR29[41] , \R_DATA_TEMPR29[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[29][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[54]  (.A(OR4_247_Y), .B(OR4_708_Y), .C(OR4_324_Y), 
        .D(OR4_650_Y), .Y(R_DATA[54]));
    OR4 OR4_30 (.A(\R_DATA_TEMPR0[60] ), .B(\R_DATA_TEMPR1[60] ), .C(
        \R_DATA_TEMPR2[60] ), .D(\R_DATA_TEMPR3[60] ), .Y(OR4_30_Y));
    OR4 OR4_650 (.A(\R_DATA_TEMPR28[54] ), .B(\R_DATA_TEMPR29[54] ), 
        .C(\R_DATA_TEMPR30[54] ), .D(\R_DATA_TEMPR31[54] ), .Y(
        OR4_650_Y));
    OR4 OR4_627 (.A(OR4_343_Y), .B(OR2_8_Y), .C(\R_DATA_TEMPR22[45] ), 
        .D(\R_DATA_TEMPR23[45] ), .Y(OR4_627_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%9%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C1 (
        .A_DOUT({\R_DATA_TEMPR9[79] , \R_DATA_TEMPR9[78] , 
        \R_DATA_TEMPR9[77] , \R_DATA_TEMPR9[76] , \R_DATA_TEMPR9[75] , 
        \R_DATA_TEMPR9[74] , \R_DATA_TEMPR9[73] , \R_DATA_TEMPR9[72] , 
        \R_DATA_TEMPR9[71] , \R_DATA_TEMPR9[70] , \R_DATA_TEMPR9[69] , 
        \R_DATA_TEMPR9[68] , \R_DATA_TEMPR9[67] , \R_DATA_TEMPR9[66] , 
        \R_DATA_TEMPR9[65] , \R_DATA_TEMPR9[64] , \R_DATA_TEMPR9[63] , 
        \R_DATA_TEMPR9[62] , \R_DATA_TEMPR9[61] , \R_DATA_TEMPR9[60] })
        , .B_DOUT({\R_DATA_TEMPR9[59] , \R_DATA_TEMPR9[58] , 
        \R_DATA_TEMPR9[57] , \R_DATA_TEMPR9[56] , \R_DATA_TEMPR9[55] , 
        \R_DATA_TEMPR9[54] , \R_DATA_TEMPR9[53] , \R_DATA_TEMPR9[52] , 
        \R_DATA_TEMPR9[51] , \R_DATA_TEMPR9[50] , \R_DATA_TEMPR9[49] , 
        \R_DATA_TEMPR9[48] , \R_DATA_TEMPR9[47] , \R_DATA_TEMPR9[46] , 
        \R_DATA_TEMPR9[45] , \R_DATA_TEMPR9[44] , \R_DATA_TEMPR9[43] , 
        \R_DATA_TEMPR9[42] , \R_DATA_TEMPR9[41] , \R_DATA_TEMPR9[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[9][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[2] , 
        \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_297 (.A(\R_DATA_TEMPR4[22] ), .B(\R_DATA_TEMPR5[22] ), .C(
        \R_DATA_TEMPR6[22] ), .D(\R_DATA_TEMPR7[22] ), .Y(OR4_297_Y));
    OR4 OR4_37 (.A(OR4_703_Y), .B(OR4_549_Y), .C(OR4_711_Y), .D(
        OR4_311_Y), .Y(OR4_37_Y));
    OR4 OR4_197 (.A(\R_DATA_TEMPR12[23] ), .B(\R_DATA_TEMPR13[23] ), 
        .C(\R_DATA_TEMPR14[23] ), .D(\R_DATA_TEMPR15[23] ), .Y(
        OR4_197_Y));
    OR4 OR4_357 (.A(\R_DATA_TEMPR16[79] ), .B(\R_DATA_TEMPR17[79] ), 
        .C(\R_DATA_TEMPR18[79] ), .D(\R_DATA_TEMPR19[79] ), .Y(
        OR4_357_Y));
    OR4 OR4_150 (.A(\R_DATA_TEMPR16[71] ), .B(\R_DATA_TEMPR17[71] ), 
        .C(\R_DATA_TEMPR18[71] ), .D(\R_DATA_TEMPR19[71] ), .Y(
        OR4_150_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[5]  (.A(CFG2_6_Y), .B(
        R_ADDR[13]), .C(R_EN), .Y(\BLKY2[5] ));
    OR4 OR4_434 (.A(OR4_679_Y), .B(OR4_541_Y), .C(OR4_528_Y), .D(
        OR4_260_Y), .Y(OR4_434_Y));
    CFG2 #( .INIT(4'h2) )  CFG2_7 (.A(W_ADDR[12]), .B(W_ADDR[11]), .Y(
        CFG2_7_Y));
    OR4 OR4_163 (.A(\R_DATA_TEMPR28[59] ), .B(\R_DATA_TEMPR29[59] ), 
        .C(\R_DATA_TEMPR30[59] ), .D(\R_DATA_TEMPR31[59] ), .Y(
        OR4_163_Y));
    OR4 OR4_343 (.A(\R_DATA_TEMPR16[45] ), .B(\R_DATA_TEMPR17[45] ), 
        .C(\R_DATA_TEMPR18[45] ), .D(\R_DATA_TEMPR19[45] ), .Y(
        OR4_343_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[7]  (.A(CFG2_5_Y), .B(
        R_ADDR[13]), .C(R_EN), .Y(\BLKY2[7] ));
    OR4 OR4_336 (.A(OR4_655_Y), .B(OR2_54_Y), .C(\R_DATA_TEMPR22[59] ), 
        .D(\R_DATA_TEMPR23[59] ), .Y(OR4_336_Y));
    OR4 OR4_415 (.A(\R_DATA_TEMPR0[31] ), .B(\R_DATA_TEMPR1[31] ), .C(
        \R_DATA_TEMPR2[31] ), .D(\R_DATA_TEMPR3[31] ), .Y(OR4_415_Y));
    OR4 OR4_442 (.A(\R_DATA_TEMPR16[51] ), .B(\R_DATA_TEMPR17[51] ), 
        .C(\R_DATA_TEMPR18[51] ), .D(\R_DATA_TEMPR19[51] ), .Y(
        OR4_442_Y));
    OR4 OR4_294 (.A(\R_DATA_TEMPR28[57] ), .B(\R_DATA_TEMPR29[57] ), 
        .C(\R_DATA_TEMPR30[57] ), .D(\R_DATA_TEMPR31[57] ), .Y(
        OR4_294_Y));
    OR4 OR4_449 (.A(\R_DATA_TEMPR12[35] ), .B(\R_DATA_TEMPR13[35] ), 
        .C(\R_DATA_TEMPR14[35] ), .D(\R_DATA_TEMPR15[35] ), .Y(
        OR4_449_Y));
    OR4 OR4_505 (.A(\R_DATA_TEMPR24[75] ), .B(\R_DATA_TEMPR25[75] ), 
        .C(\R_DATA_TEMPR26[75] ), .D(\R_DATA_TEMPR27[75] ), .Y(
        OR4_505_Y));
    OR4 \OR4_R_DATA[24]  (.A(OR4_630_Y), .B(OR4_374_Y), .C(OR4_4_Y), 
        .D(OR4_315_Y), .Y(R_DATA[24]));
    OR4 OR4_85 (.A(\R_DATA_TEMPR12[39] ), .B(\R_DATA_TEMPR13[39] ), .C(
        \R_DATA_TEMPR14[39] ), .D(\R_DATA_TEMPR15[39] ), .Y(OR4_85_Y));
    OR4 OR4_146 (.A(\R_DATA_TEMPR16[76] ), .B(\R_DATA_TEMPR17[76] ), 
        .C(\R_DATA_TEMPR18[76] ), .D(\R_DATA_TEMPR19[76] ), .Y(
        OR4_146_Y));
    OR4 OR4_158 (.A(\R_DATA_TEMPR4[57] ), .B(\R_DATA_TEMPR5[57] ), .C(
        \R_DATA_TEMPR6[57] ), .D(\R_DATA_TEMPR7[57] ), .Y(OR4_158_Y));
    OR4 \OR4_R_DATA[12]  (.A(OR4_526_Y), .B(OR4_502_Y), .C(OR4_398_Y), 
        .D(OR4_69_Y), .Y(R_DATA[12]));
    OR4 OR4_581 (.A(\R_DATA_TEMPR12[74] ), .B(\R_DATA_TEMPR13[74] ), 
        .C(\R_DATA_TEMPR14[74] ), .D(\R_DATA_TEMPR15[74] ), .Y(
        OR4_581_Y));
    OR4 OR4_575 (.A(\R_DATA_TEMPR4[5] ), .B(\R_DATA_TEMPR5[5] ), .C(
        \R_DATA_TEMPR6[5] ), .D(\R_DATA_TEMPR7[5] ), .Y(OR4_575_Y));
    OR4 \OR4_R_DATA[78]  (.A(OR4_662_Y), .B(OR4_564_Y), .C(OR4_248_Y), 
        .D(OR4_326_Y), .Y(R_DATA[78]));
    OR2 OR2_45 (.A(\R_DATA_TEMPR20[57] ), .B(\R_DATA_TEMPR21[57] ), .Y(
        OR2_45_Y));
    OR4 OR4_603 (.A(\R_DATA_TEMPR24[43] ), .B(\R_DATA_TEMPR25[43] ), 
        .C(\R_DATA_TEMPR26[43] ), .D(\R_DATA_TEMPR27[43] ), .Y(
        OR4_603_Y));
    OR4 OR4_69 (.A(\R_DATA_TEMPR28[12] ), .B(\R_DATA_TEMPR29[12] ), .C(
        \R_DATA_TEMPR30[12] ), .D(\R_DATA_TEMPR31[12] ), .Y(OR4_69_Y));
    OR2 OR2_56 (.A(\R_DATA_TEMPR20[21] ), .B(\R_DATA_TEMPR21[21] ), .Y(
        OR2_56_Y));
    OR4 OR4_227 (.A(\R_DATA_TEMPR12[73] ), .B(\R_DATA_TEMPR13[73] ), 
        .C(\R_DATA_TEMPR14[73] ), .D(\R_DATA_TEMPR15[73] ), .Y(
        OR4_227_Y));
    OR4 OR4_673 (.A(OR4_104_Y), .B(OR2_9_Y), .C(\R_DATA_TEMPR22[26] ), 
        .D(\R_DATA_TEMPR23[26] ), .Y(OR4_673_Y));
    OR4 OR4_395 (.A(\R_DATA_TEMPR24[49] ), .B(\R_DATA_TEMPR25[49] ), 
        .C(\R_DATA_TEMPR26[49] ), .D(\R_DATA_TEMPR27[49] ), .Y(
        OR4_395_Y));
    OR4 OR4_414 (.A(\R_DATA_TEMPR12[50] ), .B(\R_DATA_TEMPR13[50] ), 
        .C(\R_DATA_TEMPR14[50] ), .D(\R_DATA_TEMPR15[50] ), .Y(
        OR4_414_Y));
    OR4 OR4_127 (.A(\R_DATA_TEMPR8[65] ), .B(\R_DATA_TEMPR9[65] ), .C(
        \R_DATA_TEMPR10[65] ), .D(\R_DATA_TEMPR11[65] ), .Y(OR4_127_Y));
    OR4 OR4_348 (.A(\R_DATA_TEMPR28[74] ), .B(\R_DATA_TEMPR29[74] ), 
        .C(\R_DATA_TEMPR30[74] ), .D(\R_DATA_TEMPR31[74] ), .Y(
        OR4_348_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%30%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C1 (
        .A_DOUT({\R_DATA_TEMPR30[79] , \R_DATA_TEMPR30[78] , 
        \R_DATA_TEMPR30[77] , \R_DATA_TEMPR30[76] , 
        \R_DATA_TEMPR30[75] , \R_DATA_TEMPR30[74] , 
        \R_DATA_TEMPR30[73] , \R_DATA_TEMPR30[72] , 
        \R_DATA_TEMPR30[71] , \R_DATA_TEMPR30[70] , 
        \R_DATA_TEMPR30[69] , \R_DATA_TEMPR30[68] , 
        \R_DATA_TEMPR30[67] , \R_DATA_TEMPR30[66] , 
        \R_DATA_TEMPR30[65] , \R_DATA_TEMPR30[64] , 
        \R_DATA_TEMPR30[63] , \R_DATA_TEMPR30[62] , 
        \R_DATA_TEMPR30[61] , \R_DATA_TEMPR30[60] }), .B_DOUT({
        \R_DATA_TEMPR30[59] , \R_DATA_TEMPR30[58] , 
        \R_DATA_TEMPR30[57] , \R_DATA_TEMPR30[56] , 
        \R_DATA_TEMPR30[55] , \R_DATA_TEMPR30[54] , 
        \R_DATA_TEMPR30[53] , \R_DATA_TEMPR30[52] , 
        \R_DATA_TEMPR30[51] , \R_DATA_TEMPR30[50] , 
        \R_DATA_TEMPR30[49] , \R_DATA_TEMPR30[48] , 
        \R_DATA_TEMPR30[47] , \R_DATA_TEMPR30[46] , 
        \R_DATA_TEMPR30[45] , \R_DATA_TEMPR30[44] , 
        \R_DATA_TEMPR30[43] , \R_DATA_TEMPR30[42] , 
        \R_DATA_TEMPR30[41] , \R_DATA_TEMPR30[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[30][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_162 (.A(\R_DATA_TEMPR12[47] ), .B(\R_DATA_TEMPR13[47] ), 
        .C(\R_DATA_TEMPR14[47] ), .D(\R_DATA_TEMPR15[47] ), .Y(
        OR4_162_Y));
    OR4 OR4_282 (.A(OR4_565_Y), .B(OR4_271_Y), .C(OR4_291_Y), .D(
        OR4_663_Y), .Y(OR4_282_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%16%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0 (
        .A_DOUT({\R_DATA_TEMPR16[39] , \R_DATA_TEMPR16[38] , 
        \R_DATA_TEMPR16[37] , \R_DATA_TEMPR16[36] , 
        \R_DATA_TEMPR16[35] , \R_DATA_TEMPR16[34] , 
        \R_DATA_TEMPR16[33] , \R_DATA_TEMPR16[32] , 
        \R_DATA_TEMPR16[31] , \R_DATA_TEMPR16[30] , 
        \R_DATA_TEMPR16[29] , \R_DATA_TEMPR16[28] , 
        \R_DATA_TEMPR16[27] , \R_DATA_TEMPR16[26] , 
        \R_DATA_TEMPR16[25] , \R_DATA_TEMPR16[24] , 
        \R_DATA_TEMPR16[23] , \R_DATA_TEMPR16[22] , 
        \R_DATA_TEMPR16[21] , \R_DATA_TEMPR16[20] }), .B_DOUT({
        \R_DATA_TEMPR16[19] , \R_DATA_TEMPR16[18] , 
        \R_DATA_TEMPR16[17] , \R_DATA_TEMPR16[16] , 
        \R_DATA_TEMPR16[15] , \R_DATA_TEMPR16[14] , 
        \R_DATA_TEMPR16[13] , \R_DATA_TEMPR16[12] , 
        \R_DATA_TEMPR16[11] , \R_DATA_TEMPR16[10] , 
        \R_DATA_TEMPR16[9] , \R_DATA_TEMPR16[8] , \R_DATA_TEMPR16[7] , 
        \R_DATA_TEMPR16[6] , \R_DATA_TEMPR16[5] , \R_DATA_TEMPR16[4] , 
        \R_DATA_TEMPR16[3] , \R_DATA_TEMPR16[2] , \R_DATA_TEMPR16[1] , 
        \R_DATA_TEMPR16[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_316 (.A(OR4_379_Y), .B(OR4_53_Y), .C(OR4_328_Y), .D(
        OR4_678_Y), .Y(OR4_316_Y));
    OR2 OR2_65 (.A(\R_DATA_TEMPR20[39] ), .B(\R_DATA_TEMPR21[39] ), .Y(
        OR2_65_Y));
    OR4 OR4_134 (.A(\R_DATA_TEMPR12[69] ), .B(\R_DATA_TEMPR13[69] ), 
        .C(\R_DATA_TEMPR14[69] ), .D(\R_DATA_TEMPR15[69] ), .Y(
        OR4_134_Y));
    OR2 OR2_35 (.A(\R_DATA_TEMPR20[22] ), .B(\R_DATA_TEMPR21[22] ), .Y(
        OR2_35_Y));
    OR4 OR4_103 (.A(\R_DATA_TEMPR28[69] ), .B(\R_DATA_TEMPR29[69] ), 
        .C(\R_DATA_TEMPR30[69] ), .D(\R_DATA_TEMPR31[69] ), .Y(
        OR4_103_Y));
    OR4 OR4_224 (.A(\R_DATA_TEMPR0[3] ), .B(\R_DATA_TEMPR1[3] ), .C(
        \R_DATA_TEMPR2[3] ), .D(\R_DATA_TEMPR3[3] ), .Y(OR4_224_Y));
    OR4 OR4_149 (.A(\R_DATA_TEMPR4[8] ), .B(\R_DATA_TEMPR5[8] ), .C(
        \R_DATA_TEMPR6[8] ), .D(\R_DATA_TEMPR7[8] ), .Y(OR4_149_Y));
    OR4 OR4_380 (.A(\R_DATA_TEMPR28[14] ), .B(\R_DATA_TEMPR29[14] ), 
        .C(\R_DATA_TEMPR30[14] ), .D(\R_DATA_TEMPR31[14] ), .Y(
        OR4_380_Y));
    OR4 \OR4_R_DATA[13]  (.A(OR4_434_Y), .B(OR4_266_Y), .C(OR4_236_Y), 
        .D(OR4_219_Y), .Y(R_DATA[13]));
    OR4 OR4_173 (.A(\R_DATA_TEMPR28[16] ), .B(\R_DATA_TEMPR29[16] ), 
        .C(\R_DATA_TEMPR30[16] ), .D(\R_DATA_TEMPR31[16] ), .Y(
        OR4_173_Y));
    OR4 \OR4_R_DATA[42]  (.A(OR4_183_Y), .B(OR4_156_Y), .C(OR4_49_Y), 
        .D(OR4_448_Y), .Y(R_DATA[42]));
    OR4 OR4_269 (.A(\R_DATA_TEMPR12[75] ), .B(\R_DATA_TEMPR13[75] ), 
        .C(\R_DATA_TEMPR14[75] ), .D(\R_DATA_TEMPR15[75] ), .Y(
        OR4_269_Y));
    OR4 OR4_695 (.A(\R_DATA_TEMPR16[15] ), .B(\R_DATA_TEMPR17[15] ), 
        .C(\R_DATA_TEMPR18[15] ), .D(\R_DATA_TEMPR19[15] ), .Y(
        OR4_695_Y));
    OR4 OR4_62 (.A(OR4_216_Y), .B(OR4_625_Y), .C(OR4_51_Y), .D(
        OR4_411_Y), .Y(OR4_62_Y));
    OR4 OR4_38 (.A(OR4_377_Y), .B(OR2_37_Y), .C(\R_DATA_TEMPR22[38] ), 
        .D(\R_DATA_TEMPR23[38] ), .Y(OR4_38_Y));
    OR4 OR4_325 (.A(\R_DATA_TEMPR0[43] ), .B(\R_DATA_TEMPR1[43] ), .C(
        \R_DATA_TEMPR2[43] ), .D(\R_DATA_TEMPR3[43] ), .Y(OR4_325_Y));
    OR4 OR4_536 (.A(OR4_148_Y), .B(OR2_52_Y), .C(\R_DATA_TEMPR22[28] ), 
        .D(\R_DATA_TEMPR23[28] ), .Y(OR4_536_Y));
    OR2 OR2_50 (.A(\R_DATA_TEMPR20[60] ), .B(\R_DATA_TEMPR21[60] ), .Y(
        OR2_50_Y));
    OR4 OR4_114 (.A(\R_DATA_TEMPR4[46] ), .B(\R_DATA_TEMPR5[46] ), .C(
        \R_DATA_TEMPR6[46] ), .D(\R_DATA_TEMPR7[46] ), .Y(OR4_114_Y));
    OR4 \OR4_R_DATA[62]  (.A(OR4_19_Y), .B(OR4_716_Y), .C(OR4_618_Y), 
        .D(OR4_292_Y), .Y(R_DATA[62]));
    OR4 OR4_155 (.A(\R_DATA_TEMPR4[55] ), .B(\R_DATA_TEMPR5[55] ), .C(
        \R_DATA_TEMPR6[55] ), .D(\R_DATA_TEMPR7[55] ), .Y(OR4_155_Y));
    OR2 OR2_57 (.A(\R_DATA_TEMPR20[73] ), .B(\R_DATA_TEMPR21[73] ), .Y(
        OR2_57_Y));
    OR4 \OR4_R_DATA[79]  (.A(OR4_218_Y), .B(OR4_42_Y), .C(OR4_714_Y), 
        .D(OR4_595_Y), .Y(R_DATA[79]));
    OR4 OR4_457 (.A(\R_DATA_TEMPR24[5] ), .B(\R_DATA_TEMPR25[5] ), .C(
        \R_DATA_TEMPR26[5] ), .D(\R_DATA_TEMPR27[5] ), .Y(OR4_457_Y));
    OR4 OR4_102 (.A(\R_DATA_TEMPR16[70] ), .B(\R_DATA_TEMPR17[70] ), 
        .C(\R_DATA_TEMPR18[70] ), .D(\R_DATA_TEMPR19[70] ), .Y(
        OR4_102_Y));
    INV \INVBLKY0[0]  (.A(R_ADDR[9]), .Y(\BLKY0[0] ));
    OR4 OR4_690 (.A(OR4_91_Y), .B(OR4_527_Y), .C(OR4_675_Y), .D(
        OR4_310_Y), .Y(OR4_690_Y));
    OR4 OR4_172 (.A(\R_DATA_TEMPR12[28] ), .B(\R_DATA_TEMPR13[28] ), 
        .C(\R_DATA_TEMPR14[28] ), .D(\R_DATA_TEMPR15[28] ), .Y(
        OR4_172_Y));
    OR4 \OR4_R_DATA[51]  (.A(OR4_277_Y), .B(OR4_250_Y), .C(OR4_261_Y), 
        .D(OR4_25_Y), .Y(R_DATA[51]));
    OR4 OR4_647 (.A(\R_DATA_TEMPR24[21] ), .B(\R_DATA_TEMPR25[21] ), 
        .C(\R_DATA_TEMPR26[21] ), .D(\R_DATA_TEMPR27[21] ), .Y(
        OR4_647_Y));
    OR4 \OR4_R_DATA[43]  (.A(OR4_88_Y), .B(OR4_628_Y), .C(OR4_603_Y), 
        .D(OR4_577_Y), .Y(R_DATA[43]));
    OR4 OR4_711 (.A(\R_DATA_TEMPR8[30] ), .B(\R_DATA_TEMPR9[30] ), .C(
        \R_DATA_TEMPR10[30] ), .D(\R_DATA_TEMPR11[30] ), .Y(OR4_711_Y));
    OR4 OR4_585 (.A(\R_DATA_TEMPR12[29] ), .B(\R_DATA_TEMPR13[29] ), 
        .C(\R_DATA_TEMPR14[29] ), .D(\R_DATA_TEMPR15[29] ), .Y(
        OR4_585_Y));
    OR4 OR4_255 (.A(\R_DATA_TEMPR28[32] ), .B(\R_DATA_TEMPR29[32] ), 
        .C(\R_DATA_TEMPR30[32] ), .D(\R_DATA_TEMPR31[32] ), .Y(
        OR4_255_Y));
    OR4 OR4_397 (.A(\R_DATA_TEMPR16[17] ), .B(\R_DATA_TEMPR17[17] ), 
        .C(\R_DATA_TEMPR18[17] ), .D(\R_DATA_TEMPR19[17] ), .Y(
        OR4_397_Y));
    OR4 OR4_190 (.A(\R_DATA_TEMPR16[78] ), .B(\R_DATA_TEMPR17[78] ), 
        .C(\R_DATA_TEMPR18[78] ), .D(\R_DATA_TEMPR19[78] ), .Y(
        OR4_190_Y));
    OR4 OR4_625 (.A(\R_DATA_TEMPR4[52] ), .B(\R_DATA_TEMPR5[52] ), .C(
        \R_DATA_TEMPR6[52] ), .D(\R_DATA_TEMPR7[52] ), .Y(OR4_625_Y));
    OR4 OR4_538 (.A(\R_DATA_TEMPR8[31] ), .B(\R_DATA_TEMPR9[31] ), .C(
        \R_DATA_TEMPR10[31] ), .D(\R_DATA_TEMPR11[31] ), .Y(OR4_538_Y));
    OR4 OR4_26 (.A(\R_DATA_TEMPR28[20] ), .B(\R_DATA_TEMPR29[20] ), .C(
        \R_DATA_TEMPR30[20] ), .D(\R_DATA_TEMPR31[20] ), .Y(OR4_26_Y));
    OR4 OR4_53 (.A(\R_DATA_TEMPR4[37] ), .B(\R_DATA_TEMPR5[37] ), .C(
        \R_DATA_TEMPR6[37] ), .D(\R_DATA_TEMPR7[37] ), .Y(OR4_53_Y));
    OR4 OR4_683 (.A(\R_DATA_TEMPR0[68] ), .B(\R_DATA_TEMPR1[68] ), .C(
        \R_DATA_TEMPR2[68] ), .D(\R_DATA_TEMPR3[68] ), .Y(OR4_683_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%0%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C1 (
        .A_DOUT({\R_DATA_TEMPR0[79] , \R_DATA_TEMPR0[78] , 
        \R_DATA_TEMPR0[77] , \R_DATA_TEMPR0[76] , \R_DATA_TEMPR0[75] , 
        \R_DATA_TEMPR0[74] , \R_DATA_TEMPR0[73] , \R_DATA_TEMPR0[72] , 
        \R_DATA_TEMPR0[71] , \R_DATA_TEMPR0[70] , \R_DATA_TEMPR0[69] , 
        \R_DATA_TEMPR0[68] , \R_DATA_TEMPR0[67] , \R_DATA_TEMPR0[66] , 
        \R_DATA_TEMPR0[65] , \R_DATA_TEMPR0[64] , \R_DATA_TEMPR0[63] , 
        \R_DATA_TEMPR0[62] , \R_DATA_TEMPR0[61] , \R_DATA_TEMPR0[60] })
        , .B_DOUT({\R_DATA_TEMPR0[59] , \R_DATA_TEMPR0[58] , 
        \R_DATA_TEMPR0[57] , \R_DATA_TEMPR0[56] , \R_DATA_TEMPR0[55] , 
        \R_DATA_TEMPR0[54] , \R_DATA_TEMPR0[53] , \R_DATA_TEMPR0[52] , 
        \R_DATA_TEMPR0[51] , \R_DATA_TEMPR0[50] , \R_DATA_TEMPR0[49] , 
        \R_DATA_TEMPR0[48] , \R_DATA_TEMPR0[47] , \R_DATA_TEMPR0[46] , 
        \R_DATA_TEMPR0[45] , \R_DATA_TEMPR0[44] , \R_DATA_TEMPR0[43] , 
        \R_DATA_TEMPR0[42] , \R_DATA_TEMPR0[41] , \R_DATA_TEMPR0[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[0][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[0] , 
        \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_209 (.A(\R_DATA_TEMPR16[12] ), .B(\R_DATA_TEMPR17[12] ), 
        .C(\R_DATA_TEMPR18[12] ), .D(\R_DATA_TEMPR19[12] ), .Y(
        OR4_209_Y));
    OR4 \OR4_R_DATA[50]  (.A(OR4_131_Y), .B(OR4_300_Y), .C(OR4_632_Y), 
        .D(OR4_349_Y), .Y(R_DATA[50]));
    OR4 OR4_516 (.A(\R_DATA_TEMPR8[5] ), .B(\R_DATA_TEMPR9[5] ), .C(
        \R_DATA_TEMPR10[5] ), .D(\R_DATA_TEMPR11[5] ), .Y(OR4_516_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%15%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C1 (
        .A_DOUT({\R_DATA_TEMPR15[79] , \R_DATA_TEMPR15[78] , 
        \R_DATA_TEMPR15[77] , \R_DATA_TEMPR15[76] , 
        \R_DATA_TEMPR15[75] , \R_DATA_TEMPR15[74] , 
        \R_DATA_TEMPR15[73] , \R_DATA_TEMPR15[72] , 
        \R_DATA_TEMPR15[71] , \R_DATA_TEMPR15[70] , 
        \R_DATA_TEMPR15[69] , \R_DATA_TEMPR15[68] , 
        \R_DATA_TEMPR15[67] , \R_DATA_TEMPR15[66] , 
        \R_DATA_TEMPR15[65] , \R_DATA_TEMPR15[64] , 
        \R_DATA_TEMPR15[63] , \R_DATA_TEMPR15[62] , 
        \R_DATA_TEMPR15[61] , \R_DATA_TEMPR15[60] }), .B_DOUT({
        \R_DATA_TEMPR15[59] , \R_DATA_TEMPR15[58] , 
        \R_DATA_TEMPR15[57] , \R_DATA_TEMPR15[56] , 
        \R_DATA_TEMPR15[55] , \R_DATA_TEMPR15[54] , 
        \R_DATA_TEMPR15[53] , \R_DATA_TEMPR15[52] , 
        \R_DATA_TEMPR15[51] , \R_DATA_TEMPR15[50] , 
        \R_DATA_TEMPR15[49] , \R_DATA_TEMPR15[48] , 
        \R_DATA_TEMPR15[47] , \R_DATA_TEMPR15[46] , 
        \R_DATA_TEMPR15[45] , \R_DATA_TEMPR15[44] , 
        \R_DATA_TEMPR15[43] , \R_DATA_TEMPR15[42] , 
        \R_DATA_TEMPR15[41] , \R_DATA_TEMPR15[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[15][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%2%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0 (
        .A_DOUT({\R_DATA_TEMPR2[39] , \R_DATA_TEMPR2[38] , 
        \R_DATA_TEMPR2[37] , \R_DATA_TEMPR2[36] , \R_DATA_TEMPR2[35] , 
        \R_DATA_TEMPR2[34] , \R_DATA_TEMPR2[33] , \R_DATA_TEMPR2[32] , 
        \R_DATA_TEMPR2[31] , \R_DATA_TEMPR2[30] , \R_DATA_TEMPR2[29] , 
        \R_DATA_TEMPR2[28] , \R_DATA_TEMPR2[27] , \R_DATA_TEMPR2[26] , 
        \R_DATA_TEMPR2[25] , \R_DATA_TEMPR2[24] , \R_DATA_TEMPR2[23] , 
        \R_DATA_TEMPR2[22] , \R_DATA_TEMPR2[21] , \R_DATA_TEMPR2[20] })
        , .B_DOUT({\R_DATA_TEMPR2[19] , \R_DATA_TEMPR2[18] , 
        \R_DATA_TEMPR2[17] , \R_DATA_TEMPR2[16] , \R_DATA_TEMPR2[15] , 
        \R_DATA_TEMPR2[14] , \R_DATA_TEMPR2[13] , \R_DATA_TEMPR2[12] , 
        \R_DATA_TEMPR2[11] , \R_DATA_TEMPR2[10] , \R_DATA_TEMPR2[9] , 
        \R_DATA_TEMPR2[8] , \R_DATA_TEMPR2[7] , \R_DATA_TEMPR2[6] , 
        \R_DATA_TEMPR2[5] , \R_DATA_TEMPR2[4] , \R_DATA_TEMPR2[3] , 
        \R_DATA_TEMPR2[2] , \R_DATA_TEMPR2[1] , \R_DATA_TEMPR2[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[2][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_279 (.A(OR4_436_Y), .B(OR2_66_Y), .C(\R_DATA_TEMPR22[56] ), 
        .D(\R_DATA_TEMPR23[56] ), .Y(OR4_279_Y));
    OR4 \OR4_R_DATA[63]  (.A(OR4_658_Y), .B(OR4_469_Y), .C(OR4_435_Y), 
        .D(OR4_420_Y), .Y(R_DATA[63]));
    OR4 OR4_436 (.A(\R_DATA_TEMPR16[56] ), .B(\R_DATA_TEMPR17[56] ), 
        .C(\R_DATA_TEMPR18[56] ), .D(\R_DATA_TEMPR19[56] ), .Y(
        OR4_436_Y));
    OR4 OR4_453 (.A(\R_DATA_TEMPR4[3] ), .B(\R_DATA_TEMPR5[3] ), .C(
        \R_DATA_TEMPR6[3] ), .D(\R_DATA_TEMPR7[3] ), .Y(OR4_453_Y));
    OR4 OR4_89 (.A(\R_DATA_TEMPR16[73] ), .B(\R_DATA_TEMPR17[73] ), .C(
        \R_DATA_TEMPR18[73] ), .D(\R_DATA_TEMPR19[73] ), .Y(OR4_89_Y));
    OR4 \OR4_R_DATA[56]  (.A(OR4_608_Y), .B(OR4_279_Y), .C(OR4_401_Y), 
        .D(OR4_431_Y), .Y(R_DATA[56]));
    OR4 OR4_651 (.A(\R_DATA_TEMPR4[50] ), .B(\R_DATA_TEMPR5[50] ), .C(
        \R_DATA_TEMPR6[50] ), .D(\R_DATA_TEMPR7[50] ), .Y(OR4_651_Y));
    OR4 OR4_198 (.A(\R_DATA_TEMPR16[65] ), .B(\R_DATA_TEMPR17[65] ), 
        .C(\R_DATA_TEMPR18[65] ), .D(\R_DATA_TEMPR19[65] ), .Y(
        OR4_198_Y));
    OR4 OR4_258 (.A(OR4_587_Y), .B(OR2_16_Y), .C(\R_DATA_TEMPR22[48] ), 
        .D(\R_DATA_TEMPR23[48] ), .Y(OR4_258_Y));
    OR2 OR2_49 (.A(\R_DATA_TEMPR20[7] ), .B(\R_DATA_TEMPR21[7] ), .Y(
        OR2_49_Y));
    OR4 \OR4_R_DATA[21]  (.A(OR4_669_Y), .B(OR4_635_Y), .C(OR4_647_Y), 
        .D(OR4_416_Y), .Y(R_DATA[21]));
    OR4 OR4_620 (.A(\R_DATA_TEMPR12[43] ), .B(\R_DATA_TEMPR13[43] ), 
        .C(\R_DATA_TEMPR14[43] ), .D(\R_DATA_TEMPR15[43] ), .Y(
        OR4_620_Y));
    OR4 OR4_183 (.A(OR4_305_Y), .B(OR4_8_Y), .C(OR4_159_Y), .D(
        OR4_522_Y), .Y(OR4_183_Y));
    OR4 OR4_332 (.A(\R_DATA_TEMPR28[36] ), .B(\R_DATA_TEMPR29[36] ), 
        .C(\R_DATA_TEMPR30[36] ), .D(\R_DATA_TEMPR31[36] ), .Y(
        OR4_332_Y));
    OR4 OR4_13 (.A(\R_DATA_TEMPR28[48] ), .B(\R_DATA_TEMPR29[48] ), .C(
        \R_DATA_TEMPR30[48] ), .D(\R_DATA_TEMPR31[48] ), .Y(OR4_13_Y));
    OR4 OR4_247 (.A(OR4_106_Y), .B(OR4_276_Y), .C(OR4_346_Y), .D(
        OR4_152_Y), .Y(OR4_247_Y));
    OR4 OR4_518 (.A(\R_DATA_TEMPR16[40] ), .B(\R_DATA_TEMPR17[40] ), 
        .C(\R_DATA_TEMPR18[40] ), .D(\R_DATA_TEMPR19[40] ), .Y(
        OR4_518_Y));
    OR4 OR4_147 (.A(\R_DATA_TEMPR0[62] ), .B(\R_DATA_TEMPR1[62] ), .C(
        \R_DATA_TEMPR2[62] ), .D(\R_DATA_TEMPR3[62] ), .Y(OR4_147_Y));
    OR4 OR4_327 (.A(\R_DATA_TEMPR4[6] ), .B(\R_DATA_TEMPR5[6] ), .C(
        \R_DATA_TEMPR6[6] ), .D(\R_DATA_TEMPR7[6] ), .Y(OR4_327_Y));
    OR4 OR4_120 (.A(\R_DATA_TEMPR28[41] ), .B(\R_DATA_TEMPR29[41] ), 
        .C(\R_DATA_TEMPR30[41] ), .D(\R_DATA_TEMPR31[41] ), .Y(
        OR4_120_Y));
    OR4 OR4_51 (.A(\R_DATA_TEMPR8[52] ), .B(\R_DATA_TEMPR9[52] ), .C(
        \R_DATA_TEMPR10[52] ), .D(\R_DATA_TEMPR11[52] ), .Y(OR4_51_Y));
    INV \INVBLKY1[0]  (.A(R_ADDR[10]), .Y(\BLKY1[0] ));
    OR2 OR2_2 (.A(\R_DATA_TEMPR20[52] ), .B(\R_DATA_TEMPR21[52] ), .Y(
        OR2_2_Y));
    CFG2 #( .INIT(4'h8) )  CFG2_5 (.A(R_ADDR[12]), .B(R_ADDR[11]), .Y(
        CFG2_5_Y));
    OR4 \OR4_R_DATA[20]  (.A(OR4_534_Y), .B(OR4_698_Y), .C(OR4_301_Y), 
        .D(OR4_26_Y), .Y(R_DATA[20]));
    OR2 OR2_69 (.A(\R_DATA_TEMPR20[0] ), .B(\R_DATA_TEMPR21[0] ), .Y(
        OR2_69_Y));
    OR4 OR4_707 (.A(\R_DATA_TEMPR28[45] ), .B(\R_DATA_TEMPR29[45] ), 
        .C(\R_DATA_TEMPR30[45] ), .D(\R_DATA_TEMPR31[45] ), .Y(
        OR4_707_Y));
    OR4 OR4_704 (.A(\R_DATA_TEMPR4[29] ), .B(\R_DATA_TEMPR5[29] ), .C(
        \R_DATA_TEMPR6[29] ), .D(\R_DATA_TEMPR7[29] ), .Y(OR4_704_Y));
    OR2 OR2_39 (.A(\R_DATA_TEMPR20[31] ), .B(\R_DATA_TEMPR21[31] ), .Y(
        OR2_39_Y));
    OR4 OR4_20 (.A(\R_DATA_TEMPR8[24] ), .B(\R_DATA_TEMPR9[24] ), .C(
        \R_DATA_TEMPR10[24] ), .D(\R_DATA_TEMPR11[24] ), .Y(OR4_20_Y));
    OR4 OR4_416 (.A(\R_DATA_TEMPR28[21] ), .B(\R_DATA_TEMPR29[21] ), 
        .C(\R_DATA_TEMPR30[21] ), .D(\R_DATA_TEMPR31[21] ), .Y(
        OR4_416_Y));
    OR4 \OR4_R_DATA[26]  (.A(OR4_280_Y), .B(OR4_673_Y), .C(OR4_68_Y), 
        .D(OR4_101_Y), .Y(R_DATA[26]));
    OR4 OR4_244 (.A(\R_DATA_TEMPR12[18] ), .B(\R_DATA_TEMPR13[18] ), 
        .C(\R_DATA_TEMPR14[18] ), .D(\R_DATA_TEMPR15[18] ), .Y(
        OR4_244_Y));
    OR2 OR2_58 (.A(\R_DATA_TEMPR20[37] ), .B(\R_DATA_TEMPR21[37] ), .Y(
        OR2_58_Y));
    OR4 OR4_27 (.A(\R_DATA_TEMPR24[6] ), .B(\R_DATA_TEMPR25[6] ), .C(
        \R_DATA_TEMPR26[6] ), .D(\R_DATA_TEMPR27[6] ), .Y(OR4_27_Y));
    OR4 OR4_82 (.A(\R_DATA_TEMPR12[20] ), .B(\R_DATA_TEMPR13[20] ), .C(
        \R_DATA_TEMPR14[20] ), .D(\R_DATA_TEMPR15[20] ), .Y(OR4_82_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%15%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0 (
        .A_DOUT({\R_DATA_TEMPR15[39] , \R_DATA_TEMPR15[38] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR15[36] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR15[34] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR15[32] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR15[30] , 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR15[28] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR15[26] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR15[24] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR15[22] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR15[20] }), .B_DOUT({
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR15[18] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR15[16] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR15[14] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR15[12] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR15[10] , 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR15[8] , \R_DATA_TEMPR15[7] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR15[5] , \R_DATA_TEMPR15[4] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR15[2] , \R_DATA_TEMPR15[1] , 
        \R_DATA_TEMPR15[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_128 (.A(\R_DATA_TEMPR16[22] ), .B(\R_DATA_TEMPR17[22] ), 
        .C(\R_DATA_TEMPR18[22] ), .D(\R_DATA_TEMPR19[22] ), .Y(
        OR4_128_Y));
    OR4 OR4_230 (.A(OR4_464_Y), .B(OR4_590_Y), .C(OR4_586_Y), .D(
        OR4_710_Y), .Y(OR4_230_Y));
    OR4 OR4_537 (.A(\R_DATA_TEMPR4[68] ), .B(\R_DATA_TEMPR5[68] ), .C(
        \R_DATA_TEMPR6[68] ), .D(\R_DATA_TEMPR7[68] ), .Y(OR4_537_Y));
    OR2 OR2_42 (.A(\R_DATA_TEMPR20[8] ), .B(\R_DATA_TEMPR21[8] ), .Y(
        OR2_42_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%17%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0 (
        .A_DOUT({\R_DATA_TEMPR17[39] , \R_DATA_TEMPR17[38] , 
        \R_DATA_TEMPR17[37] , \R_DATA_TEMPR17[36] , 
        \R_DATA_TEMPR17[35] , \R_DATA_TEMPR17[34] , 
        \R_DATA_TEMPR17[33] , \R_DATA_TEMPR17[32] , 
        \R_DATA_TEMPR17[31] , \R_DATA_TEMPR17[30] , 
        \R_DATA_TEMPR17[29] , \R_DATA_TEMPR17[28] , 
        \R_DATA_TEMPR17[27] , \R_DATA_TEMPR17[26] , 
        \R_DATA_TEMPR17[25] , \R_DATA_TEMPR17[24] , 
        \R_DATA_TEMPR17[23] , \R_DATA_TEMPR17[22] , 
        \R_DATA_TEMPR17[21] , \R_DATA_TEMPR17[20] }), .B_DOUT({
        \R_DATA_TEMPR17[19] , \R_DATA_TEMPR17[18] , 
        \R_DATA_TEMPR17[17] , \R_DATA_TEMPR17[16] , 
        \R_DATA_TEMPR17[15] , \R_DATA_TEMPR17[14] , 
        \R_DATA_TEMPR17[13] , \R_DATA_TEMPR17[12] , 
        \R_DATA_TEMPR17[11] , \R_DATA_TEMPR17[10] , 
        \R_DATA_TEMPR17[9] , \R_DATA_TEMPR17[8] , \R_DATA_TEMPR17[7] , 
        \R_DATA_TEMPR17[6] , \R_DATA_TEMPR17[5] , \R_DATA_TEMPR17[4] , 
        \R_DATA_TEMPR17[3] , \R_DATA_TEMPR17[2] , \R_DATA_TEMPR17[1] , 
        \R_DATA_TEMPR17[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_182 (.A(\R_DATA_TEMPR16[16] ), .B(\R_DATA_TEMPR17[16] ), 
        .C(\R_DATA_TEMPR18[16] ), .D(\R_DATA_TEMPR19[16] ), .Y(
        OR4_182_Y));
    OR4 OR4_465 (.A(\R_DATA_TEMPR8[58] ), .B(\R_DATA_TEMPR9[58] ), .C(
        \R_DATA_TEMPR10[58] ), .D(\R_DATA_TEMPR11[58] ), .Y(OR4_465_Y));
    OR4 OR4_312 (.A(\R_DATA_TEMPR28[4] ), .B(\R_DATA_TEMPR29[4] ), .C(
        \R_DATA_TEMPR30[4] ), .D(\R_DATA_TEMPR31[4] ), .Y(OR4_312_Y));
    OR4 OR4_551 (.A(\R_DATA_TEMPR28[2] ), .B(\R_DATA_TEMPR29[2] ), .C(
        \R_DATA_TEMPR30[2] ), .D(\R_DATA_TEMPR31[2] ), .Y(OR4_551_Y));
    OR4 OR4_64 (.A(\R_DATA_TEMPR8[53] ), .B(\R_DATA_TEMPR9[53] ), .C(
        \R_DATA_TEMPR10[53] ), .D(\R_DATA_TEMPR11[53] ), .Y(OR4_64_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%23%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C1 (
        .A_DOUT({\R_DATA_TEMPR23[79] , \R_DATA_TEMPR23[78] , 
        \R_DATA_TEMPR23[77] , \R_DATA_TEMPR23[76] , 
        \R_DATA_TEMPR23[75] , \R_DATA_TEMPR23[74] , 
        \R_DATA_TEMPR23[73] , \R_DATA_TEMPR23[72] , 
        \R_DATA_TEMPR23[71] , \R_DATA_TEMPR23[70] , 
        \R_DATA_TEMPR23[69] , \R_DATA_TEMPR23[68] , 
        \R_DATA_TEMPR23[67] , \R_DATA_TEMPR23[66] , 
        \R_DATA_TEMPR23[65] , \R_DATA_TEMPR23[64] , 
        \R_DATA_TEMPR23[63] , \R_DATA_TEMPR23[62] , 
        \R_DATA_TEMPR23[61] , \R_DATA_TEMPR23[60] }), .B_DOUT({
        \R_DATA_TEMPR23[59] , \R_DATA_TEMPR23[58] , 
        \R_DATA_TEMPR23[57] , \R_DATA_TEMPR23[56] , 
        \R_DATA_TEMPR23[55] , \R_DATA_TEMPR23[54] , 
        \R_DATA_TEMPR23[53] , \R_DATA_TEMPR23[52] , 
        \R_DATA_TEMPR23[51] , \R_DATA_TEMPR23[50] , 
        \R_DATA_TEMPR23[49] , \R_DATA_TEMPR23[48] , 
        \R_DATA_TEMPR23[47] , \R_DATA_TEMPR23[46] , 
        \R_DATA_TEMPR23[45] , \R_DATA_TEMPR23[44] , 
        \R_DATA_TEMPR23[43] , \R_DATA_TEMPR23[42] , 
        \R_DATA_TEMPR23[41] , \R_DATA_TEMPR23[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[23][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[5] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_11 (.A(\R_DATA_TEMPR4[1] ), .B(\R_DATA_TEMPR5[1] ), .C(
        \R_DATA_TEMPR6[1] ), .D(\R_DATA_TEMPR7[1] ), .Y(OR4_11_Y));
    OR4 OR4_639 (.A(\R_DATA_TEMPR4[9] ), .B(\R_DATA_TEMPR5[9] ), .C(
        \R_DATA_TEMPR6[9] ), .D(\R_DATA_TEMPR7[9] ), .Y(OR4_639_Y));
    OR4 OR4_345 (.A(\R_DATA_TEMPR16[31] ), .B(\R_DATA_TEMPR17[31] ), 
        .C(\R_DATA_TEMPR18[31] ), .D(\R_DATA_TEMPR19[31] ), .Y(
        OR4_345_Y));
    OR4 OR4_236 (.A(\R_DATA_TEMPR24[13] ), .B(\R_DATA_TEMPR25[13] ), 
        .C(\R_DATA_TEMPR26[13] ), .D(\R_DATA_TEMPR27[13] ), .Y(
        OR4_236_Y));
    OR2 OR2_7 (.A(\R_DATA_TEMPR20[69] ), .B(\R_DATA_TEMPR21[69] ), .Y(
        OR2_7_Y));
    OR4 OR4_73 (.A(\R_DATA_TEMPR12[36] ), .B(\R_DATA_TEMPR13[36] ), .C(
        \R_DATA_TEMPR14[36] ), .D(\R_DATA_TEMPR15[36] ), .Y(OR4_73_Y));
    OR2 OR2_62 (.A(\R_DATA_TEMPR20[4] ), .B(\R_DATA_TEMPR21[4] ), .Y(
        OR2_62_Y));
    OR4 OR4_195 (.A(\R_DATA_TEMPR0[77] ), .B(\R_DATA_TEMPR1[77] ), .C(
        \R_DATA_TEMPR2[77] ), .D(\R_DATA_TEMPR3[77] ), .Y(OR4_195_Y));
    OR4 OR4_252 (.A(OR4_555_Y), .B(OR2_65_Y), .C(\R_DATA_TEMPR22[39] ), 
        .D(\R_DATA_TEMPR23[39] ), .Y(OR4_252_Y));
    OR4 OR4_289 (.A(\R_DATA_TEMPR4[78] ), .B(\R_DATA_TEMPR5[78] ), .C(
        \R_DATA_TEMPR6[78] ), .D(\R_DATA_TEMPR7[78] ), .Y(OR4_289_Y));
    OR4 OR4_497 (.A(OR4_61_Y), .B(OR4_304_Y), .C(OR4_619_Y), .D(
        OR4_203_Y), .Y(OR4_497_Y));
    OR2 OR2_32 (.A(\R_DATA_TEMPR20[11] ), .B(\R_DATA_TEMPR21[11] ), .Y(
        OR2_32_Y));
    OR4 OR4_634 (.A(\R_DATA_TEMPR28[58] ), .B(\R_DATA_TEMPR29[58] ), 
        .C(\R_DATA_TEMPR30[58] ), .D(\R_DATA_TEMPR31[58] ), .Y(
        OR4_634_Y));
    OR2 OR2_1 (.A(\R_DATA_TEMPR20[78] ), .B(\R_DATA_TEMPR21[78] ), .Y(
        OR2_1_Y));
    OR4 OR4_464 (.A(\R_DATA_TEMPR0[61] ), .B(\R_DATA_TEMPR1[61] ), .C(
        \R_DATA_TEMPR2[61] ), .D(\R_DATA_TEMPR3[61] ), .Y(OR4_464_Y));
    OR4 \OR4_R_DATA[57]  (.A(OR4_421_Y), .B(OR4_43_Y), .C(OR4_241_Y), 
        .D(OR4_294_Y), .Y(R_DATA[57]));
    OR4 OR4_210 (.A(\R_DATA_TEMPR24[61] ), .B(\R_DATA_TEMPR25[61] ), 
        .C(\R_DATA_TEMPR26[61] ), .D(\R_DATA_TEMPR27[61] ), .Y(
        OR4_210_Y));
    OR4 OR4_517 (.A(\R_DATA_TEMPR0[51] ), .B(\R_DATA_TEMPR1[51] ), .C(
        \R_DATA_TEMPR2[51] ), .D(\R_DATA_TEMPR3[51] ), .Y(OR4_517_Y));
    OR4 OR4_350 (.A(\R_DATA_TEMPR24[66] ), .B(\R_DATA_TEMPR25[66] ), 
        .C(\R_DATA_TEMPR26[66] ), .D(\R_DATA_TEMPR27[66] ), .Y(
        OR4_350_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%24%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0 (
        .A_DOUT({\R_DATA_TEMPR24[39] , \R_DATA_TEMPR24[38] , 
        \R_DATA_TEMPR24[37] , \R_DATA_TEMPR24[36] , 
        \R_DATA_TEMPR24[35] , \R_DATA_TEMPR24[34] , 
        \R_DATA_TEMPR24[33] , \R_DATA_TEMPR24[32] , 
        \R_DATA_TEMPR24[31] , \R_DATA_TEMPR24[30] , 
        \R_DATA_TEMPR24[29] , \R_DATA_TEMPR24[28] , 
        \R_DATA_TEMPR24[27] , \R_DATA_TEMPR24[26] , 
        \R_DATA_TEMPR24[25] , \R_DATA_TEMPR24[24] , 
        \R_DATA_TEMPR24[23] , \R_DATA_TEMPR24[22] , 
        \R_DATA_TEMPR24[21] , \R_DATA_TEMPR24[20] }), .B_DOUT({
        \R_DATA_TEMPR24[19] , \R_DATA_TEMPR24[18] , 
        \R_DATA_TEMPR24[17] , \R_DATA_TEMPR24[16] , 
        \R_DATA_TEMPR24[15] , \R_DATA_TEMPR24[14] , 
        \R_DATA_TEMPR24[13] , \R_DATA_TEMPR24[12] , 
        \R_DATA_TEMPR24[11] , \R_DATA_TEMPR24[10] , 
        \R_DATA_TEMPR24[9] , \R_DATA_TEMPR24[8] , \R_DATA_TEMPR24[7] , 
        \R_DATA_TEMPR24[6] , \R_DATA_TEMPR24[5] , \R_DATA_TEMPR24[4] , 
        \R_DATA_TEMPR24[3] , \R_DATA_TEMPR24[2] , \R_DATA_TEMPR24[1] , 
        \R_DATA_TEMPR24[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%31%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C1 (
        .A_DOUT({\R_DATA_TEMPR31[79] , \R_DATA_TEMPR31[78] , 
        \R_DATA_TEMPR31[77] , \R_DATA_TEMPR31[76] , 
        \R_DATA_TEMPR31[75] , \R_DATA_TEMPR31[74] , 
        \R_DATA_TEMPR31[73] , \R_DATA_TEMPR31[72] , 
        \R_DATA_TEMPR31[71] , \R_DATA_TEMPR31[70] , 
        \R_DATA_TEMPR31[69] , \R_DATA_TEMPR31[68] , 
        \R_DATA_TEMPR31[67] , \R_DATA_TEMPR31[66] , 
        \R_DATA_TEMPR31[65] , \R_DATA_TEMPR31[64] , 
        \R_DATA_TEMPR31[63] , \R_DATA_TEMPR31[62] , 
        \R_DATA_TEMPR31[61] , \R_DATA_TEMPR31[60] }), .B_DOUT({
        \R_DATA_TEMPR31[59] , \R_DATA_TEMPR31[58] , 
        \R_DATA_TEMPR31[57] , \R_DATA_TEMPR31[56] , 
        \R_DATA_TEMPR31[55] , \R_DATA_TEMPR31[54] , 
        \R_DATA_TEMPR31[53] , \R_DATA_TEMPR31[52] , 
        \R_DATA_TEMPR31[51] , \R_DATA_TEMPR31[50] , 
        \R_DATA_TEMPR31[49] , \R_DATA_TEMPR31[48] , 
        \R_DATA_TEMPR31[47] , \R_DATA_TEMPR31[46] , 
        \R_DATA_TEMPR31[45] , \R_DATA_TEMPR31[44] , 
        \R_DATA_TEMPR31[43] , \R_DATA_TEMPR31[42] , 
        \R_DATA_TEMPR31[41] , \R_DATA_TEMPR31[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[31][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[7] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_366 (.A(\R_DATA_TEMPR28[33] ), .B(\R_DATA_TEMPR29[33] ), 
        .C(\R_DATA_TEMPR30[33] ), .D(\R_DATA_TEMPR31[33] ), .Y(
        OR4_366_Y));
    OR4 OR4_295 (.A(\R_DATA_TEMPR8[64] ), .B(\R_DATA_TEMPR9[64] ), .C(
        \R_DATA_TEMPR10[64] ), .D(\R_DATA_TEMPR11[64] ), .Y(OR4_295_Y));
    OR4 \OR4_R_DATA[72]  (.A(OR4_495_Y), .B(OR4_476_Y), .C(OR4_372_Y), 
        .D(OR4_45_Y), .Y(R_DATA[72]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%19%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C1 (
        .A_DOUT({\R_DATA_TEMPR19[79] , \R_DATA_TEMPR19[78] , 
        \R_DATA_TEMPR19[77] , \R_DATA_TEMPR19[76] , 
        \R_DATA_TEMPR19[75] , \R_DATA_TEMPR19[74] , 
        \R_DATA_TEMPR19[73] , \R_DATA_TEMPR19[72] , 
        \R_DATA_TEMPR19[71] , \R_DATA_TEMPR19[70] , 
        \R_DATA_TEMPR19[69] , \R_DATA_TEMPR19[68] , 
        \R_DATA_TEMPR19[67] , \R_DATA_TEMPR19[66] , 
        \R_DATA_TEMPR19[65] , \R_DATA_TEMPR19[64] , 
        \R_DATA_TEMPR19[63] , \R_DATA_TEMPR19[62] , 
        \R_DATA_TEMPR19[61] , \R_DATA_TEMPR19[60] }), .B_DOUT({
        \R_DATA_TEMPR19[59] , \R_DATA_TEMPR19[58] , 
        \R_DATA_TEMPR19[57] , \R_DATA_TEMPR19[56] , 
        \R_DATA_TEMPR19[55] , \R_DATA_TEMPR19[54] , 
        \R_DATA_TEMPR19[53] , \R_DATA_TEMPR19[52] , 
        \R_DATA_TEMPR19[51] , \R_DATA_TEMPR19[50] , 
        \R_DATA_TEMPR19[49] , \R_DATA_TEMPR19[48] , 
        \R_DATA_TEMPR19[47] , \R_DATA_TEMPR19[46] , 
        \R_DATA_TEMPR19[45] , \R_DATA_TEMPR19[44] , 
        \R_DATA_TEMPR19[43] , \R_DATA_TEMPR19[42] , 
        \R_DATA_TEMPR19[41] , \R_DATA_TEMPR19[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[19][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_645 (.A(\R_DATA_TEMPR12[16] ), .B(\R_DATA_TEMPR13[16] ), 
        .C(\R_DATA_TEMPR14[16] ), .D(\R_DATA_TEMPR15[16] ), .Y(
        OR4_645_Y));
    OR4 OR4_619 (.A(\R_DATA_TEMPR8[59] ), .B(\R_DATA_TEMPR9[59] ), .C(
        \R_DATA_TEMPR10[59] ), .D(\R_DATA_TEMPR11[59] ), .Y(OR4_619_Y));
    OR4 OR4_35 (.A(\R_DATA_TEMPR4[40] ), .B(\R_DATA_TEMPR5[40] ), .C(
        \R_DATA_TEMPR6[40] ), .D(\R_DATA_TEMPR7[40] ), .Y(OR4_35_Y));
    OR4 OR4_405 (.A(\R_DATA_TEMPR0[28] ), .B(\R_DATA_TEMPR1[28] ), .C(
        \R_DATA_TEMPR2[28] ), .D(\R_DATA_TEMPR3[28] ), .Y(OR4_405_Y));
    OR4 OR4_216 (.A(\R_DATA_TEMPR0[52] ), .B(\R_DATA_TEMPR1[52] ), .C(
        \R_DATA_TEMPR2[52] ), .D(\R_DATA_TEMPR3[52] ), .Y(OR4_216_Y));
    OR4 OR4_71 (.A(\R_DATA_TEMPR8[14] ), .B(\R_DATA_TEMPR9[14] ), .C(
        \R_DATA_TEMPR10[14] ), .D(\R_DATA_TEMPR11[14] ), .Y(OR4_71_Y));
    OR4 OR4_475 (.A(\R_DATA_TEMPR0[20] ), .B(\R_DATA_TEMPR1[20] ), .C(
        \R_DATA_TEMPR2[20] ), .D(\R_DATA_TEMPR3[20] ), .Y(OR4_475_Y));
    OR4 OR4_125 (.A(OR4_638_Y), .B(OR4_488_Y), .C(OR4_365_Y), .D(
        OR4_396_Y), .Y(OR4_125_Y));
    OR4 OR4_493 (.A(\R_DATA_TEMPR24[53] ), .B(\R_DATA_TEMPR25[53] ), 
        .C(\R_DATA_TEMPR26[53] ), .D(\R_DATA_TEMPR27[53] ), .Y(
        OR4_493_Y));
    OR4 OR4_691 (.A(OR4_187_Y), .B(OR2_32_Y), .C(\R_DATA_TEMPR22[11] ), 
        .D(\R_DATA_TEMPR23[11] ), .Y(OR4_691_Y));
    OR4 OR4_614 (.A(\R_DATA_TEMPR4[17] ), .B(\R_DATA_TEMPR5[17] ), .C(
        \R_DATA_TEMPR6[17] ), .D(\R_DATA_TEMPR7[17] ), .Y(OR4_614_Y));
    OR4 OR4_427 (.A(\R_DATA_TEMPR16[1] ), .B(\R_DATA_TEMPR17[1] ), .C(
        \R_DATA_TEMPR18[1] ), .D(\R_DATA_TEMPR19[1] ), .Y(OR4_427_Y));
    OR4 OR4_298 (.A(\R_DATA_TEMPR28[75] ), .B(\R_DATA_TEMPR29[75] ), 
        .C(\R_DATA_TEMPR30[75] ), .D(\R_DATA_TEMPR31[75] ), .Y(
        OR4_298_Y));
    OR4 \OR4_R_DATA[27]  (.A(OR4_87_Y), .B(OR4_433_Y), .C(OR4_624_Y), 
        .D(OR4_692_Y), .Y(R_DATA[27]));
    OR4 OR4_28 (.A(\R_DATA_TEMPR24[65] ), .B(\R_DATA_TEMPR25[65] ), .C(
        \R_DATA_TEMPR26[65] ), .D(\R_DATA_TEMPR27[65] ), .Y(OR4_28_Y));
    OR4 OR4_640 (.A(\R_DATA_TEMPR8[51] ), .B(\R_DATA_TEMPR9[51] ), .C(
        \R_DATA_TEMPR10[51] ), .D(\R_DATA_TEMPR11[51] ), .Y(OR4_640_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%8%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0 (
        .A_DOUT({\R_DATA_TEMPR8[39] , \R_DATA_TEMPR8[38] , 
        \R_DATA_TEMPR8[37] , \R_DATA_TEMPR8[36] , \R_DATA_TEMPR8[35] , 
        \R_DATA_TEMPR8[34] , \R_DATA_TEMPR8[33] , \R_DATA_TEMPR8[32] , 
        \R_DATA_TEMPR8[31] , \R_DATA_TEMPR8[30] , \R_DATA_TEMPR8[29] , 
        \R_DATA_TEMPR8[28] , \R_DATA_TEMPR8[27] , \R_DATA_TEMPR8[26] , 
        \R_DATA_TEMPR8[25] , \R_DATA_TEMPR8[24] , \R_DATA_TEMPR8[23] , 
        \R_DATA_TEMPR8[22] , \R_DATA_TEMPR8[21] , \R_DATA_TEMPR8[20] })
        , .B_DOUT({\R_DATA_TEMPR8[19] , \R_DATA_TEMPR8[18] , 
        \R_DATA_TEMPR8[17] , \R_DATA_TEMPR8[16] , \R_DATA_TEMPR8[15] , 
        \R_DATA_TEMPR8[14] , \R_DATA_TEMPR8[13] , \R_DATA_TEMPR8[12] , 
        \R_DATA_TEMPR8[11] , \R_DATA_TEMPR8[10] , \R_DATA_TEMPR8[9] , 
        \R_DATA_TEMPR8[8] , \R_DATA_TEMPR8[7] , \R_DATA_TEMPR8[6] , 
        \R_DATA_TEMPR8[5] , \R_DATA_TEMPR8[4] , \R_DATA_TEMPR8[3] , 
        \R_DATA_TEMPR8[2] , \R_DATA_TEMPR8[1] , \R_DATA_TEMPR8[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[8][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[6]  (.A(CFG2_1_Y), .B(
        R_ADDR[13]), .C(R_EN), .Y(\BLKY2[6] ));
    OR4 \OR4_R_DATA[73]  (.A(OR4_412_Y), .B(OR4_235_Y), .C(OR4_213_Y), 
        .D(OR4_180_Y), .Y(R_DATA[73]));
    OR4 OR4_164 (.A(\R_DATA_TEMPR24[23] ), .B(\R_DATA_TEMPR25[23] ), 
        .C(\R_DATA_TEMPR26[23] ), .D(\R_DATA_TEMPR27[23] ), .Y(
        OR4_164_Y));
    OR4 OR4_404 (.A(\R_DATA_TEMPR0[65] ), .B(\R_DATA_TEMPR1[65] ), .C(
        \R_DATA_TEMPR2[65] ), .D(\R_DATA_TEMPR3[65] ), .Y(OR4_404_Y));
    OR4 OR4_225 (.A(\R_DATA_TEMPR4[4] ), .B(\R_DATA_TEMPR5[4] ), .C(
        \R_DATA_TEMPR6[4] ), .D(\R_DATA_TEMPR7[4] ), .Y(OR4_225_Y));
    CFG2 #( .INIT(4'h4) )  CFG2_2 (.A(W_ADDR[12]), .B(W_ADDR[11]), .Y(
        CFG2_2_Y));
    OR4 OR4_555 (.A(\R_DATA_TEMPR16[39] ), .B(\R_DATA_TEMPR17[39] ), 
        .C(\R_DATA_TEMPR18[39] ), .D(\R_DATA_TEMPR19[39] ), .Y(
        OR4_555_Y));
    OR4 OR4_347 (.A(\R_DATA_TEMPR8[19] ), .B(\R_DATA_TEMPR9[19] ), .C(
        \R_DATA_TEMPR10[19] ), .D(\R_DATA_TEMPR11[19] ), .Y(OR4_347_Y));
    OR4 OR4_140 (.A(\R_DATA_TEMPR16[6] ), .B(\R_DATA_TEMPR17[6] ), .C(
        \R_DATA_TEMPR18[6] ), .D(\R_DATA_TEMPR19[6] ), .Y(OR4_140_Y));
    OR4 OR4_474 (.A(\R_DATA_TEMPR0[2] ), .B(\R_DATA_TEMPR1[2] ), .C(
        \R_DATA_TEMPR2[2] ), .D(\R_DATA_TEMPR3[2] ), .Y(OR4_474_Y));
    OR4 OR4_306 (.A(\R_DATA_TEMPR16[30] ), .B(\R_DATA_TEMPR17[30] ), 
        .C(\R_DATA_TEMPR18[30] ), .D(\R_DATA_TEMPR19[30] ), .Y(
        OR4_306_Y));
    OR4 OR4_653 (.A(\R_DATA_TEMPR12[31] ), .B(\R_DATA_TEMPR13[31] ), 
        .C(\R_DATA_TEMPR14[31] ), .D(\R_DATA_TEMPR15[31] ), .Y(
        OR4_653_Y));
    CFG2 #( .INIT(4'h1) )  CFG2_3 (.A(R_ADDR[12]), .B(R_ADDR[11]), .Y(
        CFG2_3_Y));
    OR4 OR4_376 (.A(\R_DATA_TEMPR4[44] ), .B(\R_DATA_TEMPR5[44] ), .C(
        \R_DATA_TEMPR6[44] ), .D(\R_DATA_TEMPR7[44] ), .Y(OR4_376_Y));
    OR4 OR4_423 (.A(\R_DATA_TEMPR12[21] ), .B(\R_DATA_TEMPR13[21] ), 
        .C(\R_DATA_TEMPR14[21] ), .D(\R_DATA_TEMPR15[21] ), .Y(
        OR4_423_Y));
    OR4 OR4_621 (.A(\R_DATA_TEMPR28[19] ), .B(\R_DATA_TEMPR29[19] ), 
        .C(\R_DATA_TEMPR30[19] ), .D(\R_DATA_TEMPR31[19] ), .Y(
        OR4_621_Y));
    OR4 OR4_84 (.A(OR4_281_Y), .B(OR2_15_Y), .C(\R_DATA_TEMPR22[44] ), 
        .D(\R_DATA_TEMPR23[44] ), .Y(OR4_84_Y));
    OR4 OR4_148 (.A(\R_DATA_TEMPR16[28] ), .B(\R_DATA_TEMPR17[28] ), 
        .C(\R_DATA_TEMPR18[28] ), .D(\R_DATA_TEMPR19[28] ), .Y(
        OR4_148_Y));
    OR4 OR4_228 (.A(\R_DATA_TEMPR12[5] ), .B(\R_DATA_TEMPR13[5] ), .C(
        \R_DATA_TEMPR14[5] ), .D(\R_DATA_TEMPR15[5] ), .Y(OR4_228_Y));
    OR2 OR2_44 (.A(\R_DATA_TEMPR20[25] ), .B(\R_DATA_TEMPR21[25] ), .Y(
        OR2_44_Y));
    OR4 OR4_566 (.A(\R_DATA_TEMPR8[69] ), .B(\R_DATA_TEMPR9[69] ), .C(
        \R_DATA_TEMPR10[69] ), .D(\R_DATA_TEMPR11[69] ), .Y(OR4_566_Y));
    OR4 OR4_591 (.A(\R_DATA_TEMPR0[47] ), .B(\R_DATA_TEMPR1[47] ), .C(
        \R_DATA_TEMPR2[47] ), .D(\R_DATA_TEMPR3[47] ), .Y(OR4_591_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%22%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0 (
        .A_DOUT({\R_DATA_TEMPR22[39] , \R_DATA_TEMPR22[38] , 
        \R_DATA_TEMPR22[37] , \R_DATA_TEMPR22[36] , 
        \R_DATA_TEMPR22[35] , \R_DATA_TEMPR22[34] , 
        \R_DATA_TEMPR22[33] , \R_DATA_TEMPR22[32] , 
        \R_DATA_TEMPR22[31] , \R_DATA_TEMPR22[30] , 
        \R_DATA_TEMPR22[29] , \R_DATA_TEMPR22[28] , 
        \R_DATA_TEMPR22[27] , \R_DATA_TEMPR22[26] , 
        \R_DATA_TEMPR22[25] , \R_DATA_TEMPR22[24] , 
        \R_DATA_TEMPR22[23] , \R_DATA_TEMPR22[22] , 
        \R_DATA_TEMPR22[21] , \R_DATA_TEMPR22[20] }), .B_DOUT({
        \R_DATA_TEMPR22[19] , \R_DATA_TEMPR22[18] , 
        \R_DATA_TEMPR22[17] , \R_DATA_TEMPR22[16] , 
        \R_DATA_TEMPR22[15] , \R_DATA_TEMPR22[14] , 
        \R_DATA_TEMPR22[13] , \R_DATA_TEMPR22[12] , 
        \R_DATA_TEMPR22[11] , \R_DATA_TEMPR22[10] , 
        \R_DATA_TEMPR22[9] , \R_DATA_TEMPR22[8] , \R_DATA_TEMPR22[7] , 
        \R_DATA_TEMPR22[6] , \R_DATA_TEMPR22[5] , \R_DATA_TEMPR22[4] , 
        \R_DATA_TEMPR22[3] , \R_DATA_TEMPR22[2] , \R_DATA_TEMPR22[1] , 
        \R_DATA_TEMPR22[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_153 (.A(OR4_46_Y), .B(OR2_38_Y), .C(\R_DATA_TEMPR22[47] ), 
        .D(\R_DATA_TEMPR23[47] ), .Y(OR4_153_Y));
    OR4 OR4_9 (.A(OR4_319_Y), .B(OR2_79_Y), .C(\R_DATA_TEMPR22[29] ), 
        .D(\R_DATA_TEMPR23[29] ), .Y(OR4_9_Y));
    OR4 OR4_231 (.A(\R_DATA_TEMPR4[2] ), .B(\R_DATA_TEMPR5[2] ), .C(
        \R_DATA_TEMPR6[2] ), .D(\R_DATA_TEMPR7[2] ), .Y(OR4_231_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%4%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0 (
        .A_DOUT({\R_DATA_TEMPR4[39] , \R_DATA_TEMPR4[38] , 
        \R_DATA_TEMPR4[37] , \R_DATA_TEMPR4[36] , \R_DATA_TEMPR4[35] , 
        \R_DATA_TEMPR4[34] , \R_DATA_TEMPR4[33] , \R_DATA_TEMPR4[32] , 
        \R_DATA_TEMPR4[31] , \R_DATA_TEMPR4[30] , \R_DATA_TEMPR4[29] , 
        \R_DATA_TEMPR4[28] , \R_DATA_TEMPR4[27] , \R_DATA_TEMPR4[26] , 
        \R_DATA_TEMPR4[25] , \R_DATA_TEMPR4[24] , \R_DATA_TEMPR4[23] , 
        \R_DATA_TEMPR4[22] , \R_DATA_TEMPR4[21] , \R_DATA_TEMPR4[20] })
        , .B_DOUT({\R_DATA_TEMPR4[19] , \R_DATA_TEMPR4[18] , 
        \R_DATA_TEMPR4[17] , \R_DATA_TEMPR4[16] , \R_DATA_TEMPR4[15] , 
        \R_DATA_TEMPR4[14] , \R_DATA_TEMPR4[13] , \R_DATA_TEMPR4[12] , 
        \R_DATA_TEMPR4[11] , \R_DATA_TEMPR4[10] , \R_DATA_TEMPR4[9] , 
        \R_DATA_TEMPR4[8] , \R_DATA_TEMPR4[7] , \R_DATA_TEMPR4[6] , 
        \R_DATA_TEMPR4[5] , \R_DATA_TEMPR4[4] , \R_DATA_TEMPR4[3] , 
        \R_DATA_TEMPR4[2] , \R_DATA_TEMPR4[1] , \R_DATA_TEMPR4[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[4][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_104 (.A(\R_DATA_TEMPR16[26] ), .B(\R_DATA_TEMPR17[26] ), 
        .C(\R_DATA_TEMPR18[26] ), .D(\R_DATA_TEMPR19[26] ), .Y(
        OR4_104_Y));
    OR2 OR2_64 (.A(\R_DATA_TEMPR20[72] ), .B(\R_DATA_TEMPR21[72] ), .Y(
        OR2_64_Y));
    OR4 OR4_292 (.A(\R_DATA_TEMPR28[62] ), .B(\R_DATA_TEMPR29[62] ), 
        .C(\R_DATA_TEMPR30[62] ), .D(\R_DATA_TEMPR31[62] ), .Y(
        OR4_292_Y));
    OR4 OR4_174 (.A(\R_DATA_TEMPR12[6] ), .B(\R_DATA_TEMPR13[6] ), .C(
        \R_DATA_TEMPR14[6] ), .D(\R_DATA_TEMPR15[6] ), .Y(OR4_174_Y));
    OR2 OR2_34 (.A(\R_DATA_TEMPR20[63] ), .B(\R_DATA_TEMPR21[63] ), .Y(
        OR2_34_Y));
    OR4 OR4_485 (.A(\R_DATA_TEMPR8[20] ), .B(\R_DATA_TEMPR9[20] ), .C(
        \R_DATA_TEMPR10[20] ), .D(\R_DATA_TEMPR11[20] ), .Y(OR4_485_Y));
    OR4 OR4_568 (.A(\R_DATA_TEMPR4[0] ), .B(\R_DATA_TEMPR5[0] ), .C(
        \R_DATA_TEMPR6[0] ), .D(\R_DATA_TEMPR7[0] ), .Y(OR4_568_Y));
    OR4 OR4_532 (.A(\R_DATA_TEMPR24[58] ), .B(\R_DATA_TEMPR25[58] ), 
        .C(\R_DATA_TEMPR26[58] ), .D(\R_DATA_TEMPR27[58] ), .Y(
        OR4_532_Y));
    OR4 OR4_56 (.A(\R_DATA_TEMPR16[4] ), .B(\R_DATA_TEMPR17[4] ), .C(
        \R_DATA_TEMPR18[4] ), .D(\R_DATA_TEMPR19[4] ), .Y(OR4_56_Y));
    OR4 OR4_390 (.A(\R_DATA_TEMPR16[66] ), .B(\R_DATA_TEMPR17[66] ), 
        .C(\R_DATA_TEMPR18[66] ), .D(\R_DATA_TEMPR19[66] ), .Y(
        OR4_390_Y));
    OR2 OR2_55 (.A(\R_DATA_TEMPR20[19] ), .B(\R_DATA_TEMPR21[19] ), .Y(
        OR2_55_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[2]  (.A(CFG2_1_Y), .B(
        R_ADDR[13]), .C(R_EN), .Y(\BLKY2[2] ));
    OR4 OR4_701 (.A(\R_DATA_TEMPR24[35] ), .B(\R_DATA_TEMPR25[35] ), 
        .C(\R_DATA_TEMPR26[35] ), .D(\R_DATA_TEMPR27[35] ), .Y(
        OR4_701_Y));
    OR4 \OR4_R_DATA[2]  (.A(OR4_392_Y), .B(OR4_358_Y), .C(OR4_499_Y), 
        .D(OR4_551_Y), .Y(R_DATA[2]));
    OR4 OR4_521 (.A(OR4_389_Y), .B(OR2_75_Y), .C(\R_DATA_TEMPR22[53] ), 
        .D(\R_DATA_TEMPR23[53] ), .Y(OR4_521_Y));
    OR4 OR4_152 (.A(\R_DATA_TEMPR12[54] ), .B(\R_DATA_TEMPR13[54] ), 
        .C(\R_DATA_TEMPR14[54] ), .D(\R_DATA_TEMPR15[54] ), .Y(
        OR4_152_Y));
    OR4 OR4_466 (.A(\R_DATA_TEMPR8[23] ), .B(\R_DATA_TEMPR9[23] ), .C(
        \R_DATA_TEMPR10[23] ), .D(\R_DATA_TEMPR11[23] ), .Y(OR4_466_Y));
    OR4 OR4_39 (.A(\R_DATA_TEMPR24[74] ), .B(\R_DATA_TEMPR25[74] ), .C(
        \R_DATA_TEMPR26[74] ), .D(\R_DATA_TEMPR27[74] ), .Y(OR4_39_Y));
    OR4 OR4_534 (.A(OR4_475_Y), .B(OR4_317_Y), .C(OR4_485_Y), .D(
        OR4_82_Y), .Y(OR4_534_Y));
    OR4 OR4_506 (.A(\R_DATA_TEMPR0[70] ), .B(\R_DATA_TEMPR1[70] ), .C(
        \R_DATA_TEMPR2[70] ), .D(\R_DATA_TEMPR3[70] ), .Y(OR4_506_Y));
    OR4 OR4_211 (.A(\R_DATA_TEMPR16[7] ), .B(\R_DATA_TEMPR17[7] ), .C(
        \R_DATA_TEMPR18[7] ), .D(\R_DATA_TEMPR19[7] ), .Y(OR4_211_Y));
    OR4 OR4_484 (.A(\R_DATA_TEMPR0[57] ), .B(\R_DATA_TEMPR1[57] ), .C(
        \R_DATA_TEMPR2[57] ), .D(\R_DATA_TEMPR3[57] ), .Y(OR4_484_Y));
    OR2 OR2_9 (.A(\R_DATA_TEMPR20[26] ), .B(\R_DATA_TEMPR21[26] ), .Y(
        OR2_9_Y));
    OR4 OR4_576 (.A(\R_DATA_TEMPR4[62] ), .B(\R_DATA_TEMPR5[62] ), .C(
        \R_DATA_TEMPR6[62] ), .D(\R_DATA_TEMPR7[62] ), .Y(OR4_576_Y));
    OR4 OR4_145 (.A(\R_DATA_TEMPR12[10] ), .B(\R_DATA_TEMPR13[10] ), 
        .C(\R_DATA_TEMPR14[10] ), .D(\R_DATA_TEMPR15[10] ), .Y(
        OR4_145_Y));
    OR4 OR4_362 (.A(OR4_100_Y), .B(OR4_149_Y), .C(OR4_387_Y), .D(
        OR4_143_Y), .Y(OR4_362_Y));
    OR4 OR4_222 (.A(\R_DATA_TEMPR16[18] ), .B(\R_DATA_TEMPR17[18] ), 
        .C(\R_DATA_TEMPR18[18] ), .D(\R_DATA_TEMPR19[18] ), .Y(
        OR4_222_Y));
    OR4 OR4_16 (.A(\R_DATA_TEMPR12[1] ), .B(\R_DATA_TEMPR13[1] ), .C(
        \R_DATA_TEMPR14[1] ), .D(\R_DATA_TEMPR15[1] ), .Y(OR4_16_Y));
    OR4 OR4_386 (.A(\R_DATA_TEMPR16[19] ), .B(\R_DATA_TEMPR17[19] ), 
        .C(\R_DATA_TEMPR18[19] ), .D(\R_DATA_TEMPR19[19] ), .Y(
        OR4_386_Y));
    OR4 OR4_447 (.A(\R_DATA_TEMPR28[71] ), .B(\R_DATA_TEMPR29[71] ), 
        .C(\R_DATA_TEMPR30[71] ), .D(\R_DATA_TEMPR31[71] ), .Y(
        OR4_447_Y));
    OR4 OR4_259 (.A(\R_DATA_TEMPR8[34] ), .B(\R_DATA_TEMPR9[34] ), .C(
        \R_DATA_TEMPR10[34] ), .D(\R_DATA_TEMPR11[34] ), .Y(OR4_259_Y));
    OR4 OR4_4 (.A(\R_DATA_TEMPR24[24] ), .B(\R_DATA_TEMPR25[24] ), .C(
        \R_DATA_TEMPR26[24] ), .D(\R_DATA_TEMPR27[24] ), .Y(OR4_4_Y));
    OR4 OR4_331 (.A(\R_DATA_TEMPR16[27] ), .B(\R_DATA_TEMPR17[27] ), 
        .C(\R_DATA_TEMPR18[27] ), .D(\R_DATA_TEMPR19[27] ), .Y(
        OR4_331_Y));
    OR4 OR4_512 (.A(\R_DATA_TEMPR12[17] ), .B(\R_DATA_TEMPR13[17] ), 
        .C(\R_DATA_TEMPR14[17] ), .D(\R_DATA_TEMPR15[17] ), .Y(
        OR4_512_Y));
    OR4 OR4_320 (.A(\R_DATA_TEMPR28[15] ), .B(\R_DATA_TEMPR29[15] ), 
        .C(\R_DATA_TEMPR30[15] ), .D(\R_DATA_TEMPR31[15] ), .Y(
        OR4_320_Y));
    OR4 OR4_430 (.A(\R_DATA_TEMPR24[44] ), .B(\R_DATA_TEMPR25[44] ), 
        .C(\R_DATA_TEMPR26[44] ), .D(\R_DATA_TEMPR27[44] ), .Y(
        OR4_430_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%7%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0 (
        .A_DOUT({\R_DATA_TEMPR7[39] , \R_DATA_TEMPR7[38] , 
        \R_DATA_TEMPR7[37] , \R_DATA_TEMPR7[36] , \R_DATA_TEMPR7[35] , 
        \R_DATA_TEMPR7[34] , \R_DATA_TEMPR7[33] , \R_DATA_TEMPR7[32] , 
        \R_DATA_TEMPR7[31] , \R_DATA_TEMPR7[30] , \R_DATA_TEMPR7[29] , 
        \R_DATA_TEMPR7[28] , \R_DATA_TEMPR7[27] , \R_DATA_TEMPR7[26] , 
        \R_DATA_TEMPR7[25] , \R_DATA_TEMPR7[24] , \R_DATA_TEMPR7[23] , 
        \R_DATA_TEMPR7[22] , \R_DATA_TEMPR7[21] , \R_DATA_TEMPR7[20] })
        , .B_DOUT({\R_DATA_TEMPR7[19] , \R_DATA_TEMPR7[18] , 
        \R_DATA_TEMPR7[17] , \R_DATA_TEMPR7[16] , \R_DATA_TEMPR7[15] , 
        \R_DATA_TEMPR7[14] , \R_DATA_TEMPR7[13] , \R_DATA_TEMPR7[12] , 
        \R_DATA_TEMPR7[11] , \R_DATA_TEMPR7[10] , \R_DATA_TEMPR7[9] , 
        \R_DATA_TEMPR7[8] , \R_DATA_TEMPR7[7] , \R_DATA_TEMPR7[6] , 
        \R_DATA_TEMPR7[5] , \R_DATA_TEMPR7[4] , \R_DATA_TEMPR7[3] , 
        \R_DATA_TEMPR7[2] , \R_DATA_TEMPR7[1] , \R_DATA_TEMPR7[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[7][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[14]  (.A(OR4_686_Y), .B(OR4_428_Y), .C(OR4_60_Y), 
        .D(OR4_380_Y), .Y(R_DATA[14]));
    OR4 OR4_595 (.A(\R_DATA_TEMPR28[79] ), .B(\R_DATA_TEMPR29[79] ), 
        .C(\R_DATA_TEMPR30[79] ), .D(\R_DATA_TEMPR31[79] ), .Y(
        OR4_595_Y));
    OR4 OR4_245 (.A(\R_DATA_TEMPR0[56] ), .B(\R_DATA_TEMPR1[56] ), .C(
        \R_DATA_TEMPR2[56] ), .D(\R_DATA_TEMPR3[56] ), .Y(OR4_245_Y));
    OR4 OR4_508 (.A(\R_DATA_TEMPR8[12] ), .B(\R_DATA_TEMPR9[12] ), .C(
        \R_DATA_TEMPR10[12] ), .D(\R_DATA_TEMPR11[12] ), .Y(OR4_508_Y));
    OR4 OR4_50 (.A(\R_DATA_TEMPR4[35] ), .B(\R_DATA_TEMPR5[35] ), .C(
        \R_DATA_TEMPR6[35] ), .D(\R_DATA_TEMPR7[35] ), .Y(OR4_50_Y));
    OR4 OR4_514 (.A(\R_DATA_TEMPR12[53] ), .B(\R_DATA_TEMPR13[53] ), 
        .C(\R_DATA_TEMPR14[53] ), .D(\R_DATA_TEMPR15[53] ), .Y(
        OR4_514_Y));
    OR4 OR4_578 (.A(\R_DATA_TEMPR24[60] ), .B(\R_DATA_TEMPR25[60] ), 
        .C(\R_DATA_TEMPR26[60] ), .D(\R_DATA_TEMPR27[60] ), .Y(
        OR4_578_Y));
    OR4 OR4_693 (.A(\R_DATA_TEMPR8[33] ), .B(\R_DATA_TEMPR9[33] ), .C(
        \R_DATA_TEMPR10[33] ), .D(\R_DATA_TEMPR11[33] ), .Y(OR4_693_Y));
    OR4 OR4_57 (.A(\R_DATA_TEMPR16[23] ), .B(\R_DATA_TEMPR17[23] ), .C(
        \R_DATA_TEMPR18[23] ), .D(\R_DATA_TEMPR19[23] ), .Y(OR4_57_Y));
    OR4 OR4_32 (.A(\R_DATA_TEMPR28[44] ), .B(\R_DATA_TEMPR29[44] ), .C(
        \R_DATA_TEMPR30[44] ), .D(\R_DATA_TEMPR31[44] ), .Y(OR4_32_Y));
    OR4 OR4_260 (.A(\R_DATA_TEMPR12[13] ), .B(\R_DATA_TEMPR13[13] ), 
        .C(\R_DATA_TEMPR14[13] ), .D(\R_DATA_TEMPR15[13] ), .Y(
        OR4_260_Y));
    OR4 OR4_567 (.A(\R_DATA_TEMPR24[32] ), .B(\R_DATA_TEMPR25[32] ), 
        .C(\R_DATA_TEMPR26[32] ), .D(\R_DATA_TEMPR27[32] ), .Y(
        OR4_567_Y));
    OR4 OR4_406 (.A(\R_DATA_TEMPR16[50] ), .B(\R_DATA_TEMPR17[50] ), 
        .C(\R_DATA_TEMPR18[50] ), .D(\R_DATA_TEMPR19[50] ), .Y(
        OR4_406_Y));
    OR4 OR4_443 (.A(\R_DATA_TEMPR12[7] ), .B(\R_DATA_TEMPR13[7] ), .C(
        \R_DATA_TEMPR14[7] ), .D(\R_DATA_TEMPR15[7] ), .Y(OR4_443_Y));
    OR4 OR4_669 (.A(OR4_200_Y), .B(OR4_308_Y), .C(OR4_307_Y), .D(
        OR4_423_Y), .Y(OR4_669_Y));
    OR4 OR4_641 (.A(\R_DATA_TEMPR24[48] ), .B(\R_DATA_TEMPR25[48] ), 
        .C(\R_DATA_TEMPR26[48] ), .D(\R_DATA_TEMPR27[48] ), .Y(
        OR4_641_Y));
    OR4 OR4_476 (.A(OR4_165_Y), .B(OR2_64_Y), .C(\R_DATA_TEMPR22[72] ), 
        .D(\R_DATA_TEMPR23[72] ), .Y(OR4_476_Y));
    OR4 OR4_184 (.A(\R_DATA_TEMPR0[63] ), .B(\R_DATA_TEMPR1[63] ), .C(
        \R_DATA_TEMPR2[63] ), .D(\R_DATA_TEMPR3[63] ), .Y(OR4_184_Y));
    OR4 OR4_311 (.A(\R_DATA_TEMPR12[30] ), .B(\R_DATA_TEMPR13[30] ), 
        .C(\R_DATA_TEMPR14[30] ), .D(\R_DATA_TEMPR15[30] ), .Y(
        OR4_311_Y));
    OR4 OR4_248 (.A(\R_DATA_TEMPR24[78] ), .B(\R_DATA_TEMPR25[78] ), 
        .C(\R_DATA_TEMPR26[78] ), .D(\R_DATA_TEMPR27[78] ), .Y(
        OR4_248_Y));
    OR4 OR4_302 (.A(\R_DATA_TEMPR24[36] ), .B(\R_DATA_TEMPR25[36] ), 
        .C(\R_DATA_TEMPR26[36] ), .D(\R_DATA_TEMPR27[36] ), .Y(
        OR4_302_Y));
    OR4 OR4_266 (.A(OR4_113_Y), .B(OR2_76_Y), .C(\R_DATA_TEMPR22[13] ), 
        .D(\R_DATA_TEMPR23[13] ), .Y(OR4_266_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%8%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C1 (
        .A_DOUT({\R_DATA_TEMPR8[79] , \R_DATA_TEMPR8[78] , 
        \R_DATA_TEMPR8[77] , \R_DATA_TEMPR8[76] , \R_DATA_TEMPR8[75] , 
        \R_DATA_TEMPR8[74] , \R_DATA_TEMPR8[73] , \R_DATA_TEMPR8[72] , 
        \R_DATA_TEMPR8[71] , \R_DATA_TEMPR8[70] , \R_DATA_TEMPR8[69] , 
        \R_DATA_TEMPR8[68] , \R_DATA_TEMPR8[67] , \R_DATA_TEMPR8[66] , 
        \R_DATA_TEMPR8[65] , \R_DATA_TEMPR8[64] , \R_DATA_TEMPR8[63] , 
        \R_DATA_TEMPR8[62] , \R_DATA_TEMPR8[61] , \R_DATA_TEMPR8[60] })
        , .B_DOUT({\R_DATA_TEMPR8[59] , \R_DATA_TEMPR8[58] , 
        \R_DATA_TEMPR8[57] , \R_DATA_TEMPR8[56] , \R_DATA_TEMPR8[55] , 
        \R_DATA_TEMPR8[54] , \R_DATA_TEMPR8[53] , \R_DATA_TEMPR8[52] , 
        \R_DATA_TEMPR8[51] , \R_DATA_TEMPR8[50] , \R_DATA_TEMPR8[49] , 
        \R_DATA_TEMPR8[48] , \R_DATA_TEMPR8[47] , \R_DATA_TEMPR8[46] , 
        \R_DATA_TEMPR8[45] , \R_DATA_TEMPR8[44] , \R_DATA_TEMPR8[43] , 
        \R_DATA_TEMPR8[42] , \R_DATA_TEMPR8[41] , \R_DATA_TEMPR8[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[8][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[2] , 
        \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_10 (.A(\R_DATA_TEMPR24[40] ), .B(\R_DATA_TEMPR25[40] ), .C(
        \R_DATA_TEMPR26[40] ), .D(\R_DATA_TEMPR27[40] ), .Y(OR4_10_Y));
    OR4 OR4_25 (.A(\R_DATA_TEMPR28[51] ), .B(\R_DATA_TEMPR29[51] ), .C(
        \R_DATA_TEMPR30[51] ), .D(\R_DATA_TEMPR31[51] ), .Y(OR4_25_Y));
    OR4 OR4_76 (.A(\R_DATA_TEMPR28[10] ), .B(\R_DATA_TEMPR29[10] ), .C(
        \R_DATA_TEMPR30[10] ), .D(\R_DATA_TEMPR31[10] ), .Y(OR4_76_Y));
    OR4 OR4_410 (.A(\R_DATA_TEMPR4[49] ), .B(\R_DATA_TEMPR5[49] ), .C(
        \R_DATA_TEMPR6[49] ), .D(\R_DATA_TEMPR7[49] ), .Y(OR4_410_Y));
    OR4 OR4_339 (.A(\R_DATA_TEMPR24[22] ), .B(\R_DATA_TEMPR25[22] ), 
        .C(\R_DATA_TEMPR26[22] ), .D(\R_DATA_TEMPR27[22] ), .Y(
        OR4_339_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[4]  (.A(CFG2_4_Y), .B(
        W_ADDR[13]), .C(W_EN), .Y(\BLKX2[4] ));
    OR4 OR4_193 (.A(OR4_394_Y), .B(OR2_63_Y), .C(\R_DATA_TEMPR22[61] ), 
        .D(\R_DATA_TEMPR23[61] ), .Y(OR4_193_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%4%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C1 (
        .A_DOUT({\R_DATA_TEMPR4[79] , \R_DATA_TEMPR4[78] , 
        \R_DATA_TEMPR4[77] , \R_DATA_TEMPR4[76] , \R_DATA_TEMPR4[75] , 
        \R_DATA_TEMPR4[74] , \R_DATA_TEMPR4[73] , \R_DATA_TEMPR4[72] , 
        \R_DATA_TEMPR4[71] , \R_DATA_TEMPR4[70] , \R_DATA_TEMPR4[69] , 
        \R_DATA_TEMPR4[68] , \R_DATA_TEMPR4[67] , \R_DATA_TEMPR4[66] , 
        \R_DATA_TEMPR4[65] , \R_DATA_TEMPR4[64] , \R_DATA_TEMPR4[63] , 
        \R_DATA_TEMPR4[62] , \R_DATA_TEMPR4[61] , \R_DATA_TEMPR4[60] })
        , .B_DOUT({\R_DATA_TEMPR4[59] , \R_DATA_TEMPR4[58] , 
        \R_DATA_TEMPR4[57] , \R_DATA_TEMPR4[56] , \R_DATA_TEMPR4[55] , 
        \R_DATA_TEMPR4[54] , \R_DATA_TEMPR4[53] , \R_DATA_TEMPR4[52] , 
        \R_DATA_TEMPR4[51] , \R_DATA_TEMPR4[50] , \R_DATA_TEMPR4[49] , 
        \R_DATA_TEMPR4[48] , \R_DATA_TEMPR4[47] , \R_DATA_TEMPR4[46] , 
        \R_DATA_TEMPR4[45] , \R_DATA_TEMPR4[44] , \R_DATA_TEMPR4[43] , 
        \R_DATA_TEMPR4[42] , \R_DATA_TEMPR4[41] , \R_DATA_TEMPR4[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[4][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[1] , 
        \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_372 (.A(\R_DATA_TEMPR24[72] ), .B(\R_DATA_TEMPR25[72] ), 
        .C(\R_DATA_TEMPR26[72] ), .D(\R_DATA_TEMPR27[72] ), .Y(
        OR4_372_Y));
    OR4 \OR4_R_DATA[44]  (.A(OR4_335_Y), .B(OR4_84_Y), .C(OR4_430_Y), 
        .D(OR4_32_Y), .Y(R_DATA[44]));
    OR4 OR4_525 (.A(\R_DATA_TEMPR8[0] ), .B(\R_DATA_TEMPR9[0] ), .C(
        \R_DATA_TEMPR10[0] ), .D(\R_DATA_TEMPR11[0] ), .Y(OR4_525_Y));
    OR4 OR4_17 (.A(\R_DATA_TEMPR4[56] ), .B(\R_DATA_TEMPR5[56] ), .C(
        \R_DATA_TEMPR6[56] ), .D(\R_DATA_TEMPR7[56] ), .Y(OR4_17_Y));
    OR4 OR4_664 (.A(OR4_150_Y), .B(OR2_3_Y), .C(\R_DATA_TEMPR22[71] ), 
        .D(\R_DATA_TEMPR23[71] ), .Y(OR4_664_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%13%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C1 (
        .A_DOUT({\R_DATA_TEMPR13[79] , \R_DATA_TEMPR13[78] , 
        \R_DATA_TEMPR13[77] , \R_DATA_TEMPR13[76] , 
        \R_DATA_TEMPR13[75] , \R_DATA_TEMPR13[74] , 
        \R_DATA_TEMPR13[73] , \R_DATA_TEMPR13[72] , 
        \R_DATA_TEMPR13[71] , \R_DATA_TEMPR13[70] , 
        \R_DATA_TEMPR13[69] , \R_DATA_TEMPR13[68] , 
        \R_DATA_TEMPR13[67] , \R_DATA_TEMPR13[66] , 
        \R_DATA_TEMPR13[65] , \R_DATA_TEMPR13[64] , 
        \R_DATA_TEMPR13[63] , \R_DATA_TEMPR13[62] , 
        \R_DATA_TEMPR13[61] , \R_DATA_TEMPR13[60] }), .B_DOUT({
        \R_DATA_TEMPR13[59] , \R_DATA_TEMPR13[58] , 
        \R_DATA_TEMPR13[57] , \R_DATA_TEMPR13[56] , 
        \R_DATA_TEMPR13[55] , \R_DATA_TEMPR13[54] , 
        \R_DATA_TEMPR13[53] , \R_DATA_TEMPR13[52] , 
        \R_DATA_TEMPR13[51] , \R_DATA_TEMPR13[50] , 
        \R_DATA_TEMPR13[49] , \R_DATA_TEMPR13[48] , 
        \R_DATA_TEMPR13[47] , \R_DATA_TEMPR13[46] , 
        \R_DATA_TEMPR13[45] , \R_DATA_TEMPR13[44] , 
        \R_DATA_TEMPR13[43] , \R_DATA_TEMPR13[42] , 
        \R_DATA_TEMPR13[41] , \R_DATA_TEMPR13[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[13][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_623 (.A(\R_DATA_TEMPR0[41] ), .B(\R_DATA_TEMPR1[41] ), .C(
        \R_DATA_TEMPR2[41] ), .D(\R_DATA_TEMPR3[41] ), .Y(OR4_623_Y));
    OR4 OR4_586 (.A(\R_DATA_TEMPR8[61] ), .B(\R_DATA_TEMPR9[61] ), .C(
        \R_DATA_TEMPR10[61] ), .D(\R_DATA_TEMPR11[61] ), .Y(OR4_586_Y));
    OR4 OR4_200 (.A(\R_DATA_TEMPR0[21] ), .B(\R_DATA_TEMPR1[21] ), .C(
        \R_DATA_TEMPR2[21] ), .D(\R_DATA_TEMPR3[21] ), .Y(OR4_200_Y));
    OR4 \OR4_R_DATA[64]  (.A(OR4_189_Y), .B(OR4_652_Y), .C(OR4_283_Y), 
        .D(OR4_598_Y), .Y(R_DATA[64]));
    OR4 OR4_507 (.A(\R_DATA_TEMPR4[73] ), .B(\R_DATA_TEMPR5[73] ), .C(
        \R_DATA_TEMPR6[73] ), .D(\R_DATA_TEMPR7[73] ), .Y(OR4_507_Y));
    OR2 OR2_59 (.A(\R_DATA_TEMPR20[46] ), .B(\R_DATA_TEMPR21[46] ), .Y(
        OR2_59_Y));
    OR4 OR4_270 (.A(\R_DATA_TEMPR12[44] ), .B(\R_DATA_TEMPR13[44] ), 
        .C(\R_DATA_TEMPR14[44] ), .D(\R_DATA_TEMPR15[44] ), .Y(
        OR4_270_Y));
    OR4 OR4_577 (.A(\R_DATA_TEMPR28[43] ), .B(\R_DATA_TEMPR29[43] ), 
        .C(\R_DATA_TEMPR30[43] ), .D(\R_DATA_TEMPR31[43] ), .Y(
        OR4_577_Y));
    OR4 OR4_541 (.A(\R_DATA_TEMPR4[13] ), .B(\R_DATA_TEMPR5[13] ), .C(
        \R_DATA_TEMPR6[13] ), .D(\R_DATA_TEMPR7[13] ), .Y(OR4_541_Y));
    OR4 OR4_192 (.A(\R_DATA_TEMPR12[56] ), .B(\R_DATA_TEMPR13[56] ), 
        .C(\R_DATA_TEMPR14[56] ), .D(\R_DATA_TEMPR15[56] ), .Y(
        OR4_192_Y));
    OR4 OR4_319 (.A(\R_DATA_TEMPR16[29] ), .B(\R_DATA_TEMPR17[29] ), 
        .C(\R_DATA_TEMPR18[29] ), .D(\R_DATA_TEMPR19[29] ), .Y(
        OR4_319_Y));
    OR4 OR4_609 (.A(\R_DATA_TEMPR12[48] ), .B(\R_DATA_TEMPR13[48] ), 
        .C(\R_DATA_TEMPR14[48] ), .D(\R_DATA_TEMPR15[48] ), .Y(
        OR4_609_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%28%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C1 (
        .A_DOUT({\R_DATA_TEMPR28[79] , \R_DATA_TEMPR28[78] , 
        \R_DATA_TEMPR28[77] , \R_DATA_TEMPR28[76] , 
        \R_DATA_TEMPR28[75] , \R_DATA_TEMPR28[74] , 
        \R_DATA_TEMPR28[73] , \R_DATA_TEMPR28[72] , 
        \R_DATA_TEMPR28[71] , \R_DATA_TEMPR28[70] , 
        \R_DATA_TEMPR28[69] , \R_DATA_TEMPR28[68] , 
        \R_DATA_TEMPR28[67] , \R_DATA_TEMPR28[66] , 
        \R_DATA_TEMPR28[65] , \R_DATA_TEMPR28[64] , 
        \R_DATA_TEMPR28[63] , \R_DATA_TEMPR28[62] , 
        \R_DATA_TEMPR28[61] , \R_DATA_TEMPR28[60] }), .B_DOUT({
        \R_DATA_TEMPR28[59] , \R_DATA_TEMPR28[58] , 
        \R_DATA_TEMPR28[57] , \R_DATA_TEMPR28[56] , 
        \R_DATA_TEMPR28[55] , \R_DATA_TEMPR28[54] , 
        \R_DATA_TEMPR28[53] , \R_DATA_TEMPR28[52] , 
        \R_DATA_TEMPR28[51] , \R_DATA_TEMPR28[50] , 
        \R_DATA_TEMPR28[49] , \R_DATA_TEMPR28[48] , 
        \R_DATA_TEMPR28[47] , \R_DATA_TEMPR28[46] , 
        \R_DATA_TEMPR28[45] , \R_DATA_TEMPR28[44] , 
        \R_DATA_TEMPR28[43] , \R_DATA_TEMPR28[42] , 
        \R_DATA_TEMPR28[41] , \R_DATA_TEMPR28[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[28][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_123 (.A(\R_DATA_TEMPR0[25] ), .B(\R_DATA_TEMPR1[25] ), .C(
        \R_DATA_TEMPR2[25] ), .D(\R_DATA_TEMPR3[25] ), .Y(OR4_123_Y));
    OR4 OR4_679 (.A(\R_DATA_TEMPR0[13] ), .B(\R_DATA_TEMPR1[13] ), .C(
        \R_DATA_TEMPR2[13] ), .D(\R_DATA_TEMPR3[13] ), .Y(OR4_679_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%14%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0 (
        .A_DOUT({\R_DATA_TEMPR14[39] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR14[37] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR14[35] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR14[33] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR14[31] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR14[29] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR14[27] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR14[25] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR14[23] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR14[21] , \R_DATA_TEMPR14[20] }), .B_DOUT({
        \R_DATA_TEMPR14[19] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR14[17] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR14[15] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR14[13] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR14[11] , \R_DATA_TEMPR14[10] , 
        \R_DATA_TEMPR14[9] , \R_DATA_TEMPR14[8] , \R_DATA_TEMPR14[7] , 
        \R_DATA_TEMPR14[6] , \R_DATA_TEMPR14[5] , \R_DATA_TEMPR14[4] , 
        \R_DATA_TEMPR14[3] , \R_DATA_TEMPR14[2] , \R_DATA_TEMPR14[1] , 
        \R_DATA_TEMPR14[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_206 (.A(OR4_57_Y), .B(OR2_24_Y), .C(\R_DATA_TEMPR22[23] ), 
        .D(\R_DATA_TEMPR23[23] ), .Y(OR4_206_Y));
    OR4 OR4_533 (.A(\R_DATA_TEMPR8[7] ), .B(\R_DATA_TEMPR9[7] ), .C(
        \R_DATA_TEMPR10[7] ), .D(\R_DATA_TEMPR11[7] ), .Y(OR4_533_Y));
    CFG2 #( .INIT(4'h2) )  CFG2_1 (.A(R_ADDR[12]), .B(R_ADDR[11]), .Y(
        CFG2_1_Y));
    OR4 OR4_70 (.A(\R_DATA_TEMPR24[55] ), .B(\R_DATA_TEMPR25[55] ), .C(
        \R_DATA_TEMPR26[55] ), .D(\R_DATA_TEMPR27[55] ), .Y(OR4_70_Y));
    OR4 OR4_588 (.A(\R_DATA_TEMPR4[58] ), .B(\R_DATA_TEMPR5[58] ), .C(
        \R_DATA_TEMPR6[58] ), .D(\R_DATA_TEMPR7[58] ), .Y(OR4_588_Y));
    OR4 OR4_58 (.A(\R_DATA_TEMPR28[39] ), .B(\R_DATA_TEMPR29[39] ), .C(
        \R_DATA_TEMPR30[39] ), .D(\R_DATA_TEMPR31[39] ), .Y(OR4_58_Y));
    OR4 OR4_276 (.A(\R_DATA_TEMPR4[54] ), .B(\R_DATA_TEMPR5[54] ), .C(
        \R_DATA_TEMPR6[54] ), .D(\R_DATA_TEMPR7[54] ), .Y(OR4_276_Y));
    OR4 OR4_242 (.A(OR4_375_Y), .B(OR2_10_Y), .C(\R_DATA_TEMPR22[9] ), 
        .D(\R_DATA_TEMPR23[9] ), .Y(OR4_242_Y));
    OR4 OR4_77 (.A(\R_DATA_TEMPR8[35] ), .B(\R_DATA_TEMPR9[35] ), .C(
        \R_DATA_TEMPR10[35] ), .D(\R_DATA_TEMPR11[35] ), .Y(OR4_77_Y));
    OR4 OR4_604 (.A(OR4_65_Y), .B(OR2_36_Y), .C(\R_DATA_TEMPR22[34] ), 
        .D(\R_DATA_TEMPR23[34] ), .Y(OR4_604_Y));
    OR4 OR4_299 (.A(\R_DATA_TEMPR28[60] ), .B(\R_DATA_TEMPR29[60] ), 
        .C(\R_DATA_TEMPR30[60] ), .D(\R_DATA_TEMPR31[60] ), .Y(
        OR4_299_Y));
    OR4 OR4_674 (.A(\R_DATA_TEMPR24[71] ), .B(\R_DATA_TEMPR25[71] ), 
        .C(\R_DATA_TEMPR26[71] ), .D(\R_DATA_TEMPR27[71] ), .Y(
        OR4_674_Y));
    OR4 OR4_455 (.A(\R_DATA_TEMPR12[71] ), .B(\R_DATA_TEMPR13[71] ), 
        .C(\R_DATA_TEMPR14[71] ), .D(\R_DATA_TEMPR15[71] ), .Y(
        OR4_455_Y));
    OR4 OR4_486 (.A(\R_DATA_TEMPR8[72] ), .B(\R_DATA_TEMPR9[72] ), .C(
        \R_DATA_TEMPR10[72] ), .D(\R_DATA_TEMPR11[72] ), .Y(OR4_486_Y));
    OR4 \OR4_R_DATA[5]  (.A(OR4_107_Y), .B(OR4_688_Y), .C(OR4_457_Y), 
        .D(OR4_601_Y), .Y(R_DATA[5]));
    OR2 OR2_52 (.A(\R_DATA_TEMPR20[28] ), .B(\R_DATA_TEMPR21[28] ), .Y(
        OR2_52_Y));
    OR4 OR4_340 (.A(\R_DATA_TEMPR16[36] ), .B(\R_DATA_TEMPR17[36] ), 
        .C(\R_DATA_TEMPR18[36] ), .D(\R_DATA_TEMPR19[36] ), .Y(
        OR4_340_Y));
    OR4 OR4_719 (.A(\R_DATA_TEMPR8[49] ), .B(\R_DATA_TEMPR9[49] ), .C(
        \R_DATA_TEMPR10[49] ), .D(\R_DATA_TEMPR11[49] ), .Y(OR4_719_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%26%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C1 (
        .A_DOUT({\R_DATA_TEMPR26[79] , \R_DATA_TEMPR26[78] , 
        \R_DATA_TEMPR26[77] , \R_DATA_TEMPR26[76] , 
        \R_DATA_TEMPR26[75] , \R_DATA_TEMPR26[74] , 
        \R_DATA_TEMPR26[73] , \R_DATA_TEMPR26[72] , 
        \R_DATA_TEMPR26[71] , \R_DATA_TEMPR26[70] , 
        \R_DATA_TEMPR26[69] , \R_DATA_TEMPR26[68] , 
        \R_DATA_TEMPR26[67] , \R_DATA_TEMPR26[66] , 
        \R_DATA_TEMPR26[65] , \R_DATA_TEMPR26[64] , 
        \R_DATA_TEMPR26[63] , \R_DATA_TEMPR26[62] , 
        \R_DATA_TEMPR26[61] , \R_DATA_TEMPR26[60] }), .B_DOUT({
        \R_DATA_TEMPR26[59] , \R_DATA_TEMPR26[58] , 
        \R_DATA_TEMPR26[57] , \R_DATA_TEMPR26[56] , 
        \R_DATA_TEMPR26[55] , \R_DATA_TEMPR26[54] , 
        \R_DATA_TEMPR26[53] , \R_DATA_TEMPR26[52] , 
        \R_DATA_TEMPR26[51] , \R_DATA_TEMPR26[50] , 
        \R_DATA_TEMPR26[49] , \R_DATA_TEMPR26[48] , 
        \R_DATA_TEMPR26[47] , \R_DATA_TEMPR26[46] , 
        \R_DATA_TEMPR26[45] , \R_DATA_TEMPR26[44] , 
        \R_DATA_TEMPR26[43] , \R_DATA_TEMPR26[42] , 
        \R_DATA_TEMPR26[41] , \R_DATA_TEMPR26[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[26][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[11]  (.A(OR4_2_Y), .B(OR4_691_Y), .C(OR4_706_Y), 
        .D(OR4_481_Y), .Y(R_DATA[11]));
    OR4 OR4_122 (.A(OR4_14_Y), .B(OR4_166_Y), .C(OR4_259_Y), .D(
        OR4_47_Y), .Y(OR4_122_Y));
    OR4 OR4_382 (.A(\R_DATA_TEMPR4[10] ), .B(\R_DATA_TEMPR5[10] ), .C(
        \R_DATA_TEMPR6[10] ), .D(\R_DATA_TEMPR7[10] ), .Y(OR4_382_Y));
    OR4 \OR4_R_DATA[9]  (.A(OR4_90_Y), .B(OR4_242_Y), .C(OR4_417_Y), 
        .D(OR4_560_Y), .Y(R_DATA[9]));
    OR4 OR4_18 (.A(\R_DATA_TEMPR28[22] ), .B(\R_DATA_TEMPR29[22] ), .C(
        \R_DATA_TEMPR30[22] ), .D(\R_DATA_TEMPR31[22] ), .Y(OR4_18_Y));
    OR4 OR4_513 (.A(\R_DATA_TEMPR8[70] ), .B(\R_DATA_TEMPR9[70] ), .C(
        \R_DATA_TEMPR10[70] ), .D(\R_DATA_TEMPR11[70] ), .Y(OR4_513_Y));
    OR4 OR4_34 (.A(OR4_138_Y), .B(OR2_12_Y), .C(\R_DATA_TEMPR22[10] ), 
        .D(\R_DATA_TEMPR23[10] ), .Y(OR4_34_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%0%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0 (
        .A_DOUT({\R_DATA_TEMPR0[39] , \R_DATA_TEMPR0[38] , 
        \R_DATA_TEMPR0[37] , \R_DATA_TEMPR0[36] , \R_DATA_TEMPR0[35] , 
        \R_DATA_TEMPR0[34] , \R_DATA_TEMPR0[33] , \R_DATA_TEMPR0[32] , 
        \R_DATA_TEMPR0[31] , \R_DATA_TEMPR0[30] , \R_DATA_TEMPR0[29] , 
        \R_DATA_TEMPR0[28] , \R_DATA_TEMPR0[27] , \R_DATA_TEMPR0[26] , 
        \R_DATA_TEMPR0[25] , \R_DATA_TEMPR0[24] , \R_DATA_TEMPR0[23] , 
        \R_DATA_TEMPR0[22] , \R_DATA_TEMPR0[21] , \R_DATA_TEMPR0[20] })
        , .B_DOUT({\R_DATA_TEMPR0[19] , \R_DATA_TEMPR0[18] , 
        \R_DATA_TEMPR0[17] , \R_DATA_TEMPR0[16] , \R_DATA_TEMPR0[15] , 
        \R_DATA_TEMPR0[14] , \R_DATA_TEMPR0[13] , \R_DATA_TEMPR0[12] , 
        \R_DATA_TEMPR0[11] , \R_DATA_TEMPR0[10] , \R_DATA_TEMPR0[9] , 
        \R_DATA_TEMPR0[8] , \R_DATA_TEMPR0[7] , \R_DATA_TEMPR0[6] , 
        \R_DATA_TEMPR0[5] , \R_DATA_TEMPR0[4] , \R_DATA_TEMPR0[3] , 
        \R_DATA_TEMPR0[2] , \R_DATA_TEMPR0[1] , \R_DATA_TEMPR0[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[0][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_454 (.A(\R_DATA_TEMPR28[40] ), .B(\R_DATA_TEMPR29[40] ), 
        .C(\R_DATA_TEMPR30[40] ), .D(\R_DATA_TEMPR31[40] ), .Y(
        OR4_454_Y));
    OR4 \OR4_R_DATA[35]  (.A(OR4_67_Y), .B(OR4_418_Y), .C(OR4_701_Y), 
        .D(OR4_494_Y), .Y(R_DATA[35]));
    OR4 \OR4_R_DATA[10]  (.A(OR4_593_Y), .B(OR4_34_Y), .C(OR4_359_Y), 
        .D(OR4_76_Y), .Y(R_DATA[10]));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[1]  (.A(CFG2_2_Y), .B(
        W_ADDR[13]), .C(W_EN), .Y(\BLKX2[1] ));
    OR4 OR4_229 (.A(\R_DATA_TEMPR0[71] ), .B(\R_DATA_TEMPR1[71] ), .C(
        \R_DATA_TEMPR2[71] ), .D(\R_DATA_TEMPR3[71] ), .Y(OR4_229_Y));
    OR4 OR4_356 (.A(\R_DATA_TEMPR4[12] ), .B(\R_DATA_TEMPR5[12] ), .C(
        \R_DATA_TEMPR6[12] ), .D(\R_DATA_TEMPR7[12] ), .Y(OR4_356_Y));
    OR4 OR4_261 (.A(\R_DATA_TEMPR24[51] ), .B(\R_DATA_TEMPR25[51] ), 
        .C(\R_DATA_TEMPR26[51] ), .D(\R_DATA_TEMPR27[51] ), .Y(
        OR4_261_Y));
    OR2 OR2_23 (.A(\R_DATA_TEMPR20[77] ), .B(\R_DATA_TEMPR21[77] ), .Y(
        OR2_23_Y));
    OR4 OR4_29 (.A(\R_DATA_TEMPR28[17] ), .B(\R_DATA_TEMPR29[17] ), .C(
        \R_DATA_TEMPR30[17] ), .D(\R_DATA_TEMPR31[17] ), .Y(OR4_29_Y));
    OR4 \OR4_R_DATA[16]  (.A(OR4_330_Y), .B(OR4_6_Y), .C(OR4_129_Y), 
        .D(OR4_173_Y), .Y(R_DATA[16]));
    OR4 OR4_280 (.A(OR4_629_Y), .B(OR4_407_Y), .C(OR4_446_Y), .D(
        OR4_579_Y), .Y(OR4_280_Y));
    OR4 OR4_587 (.A(\R_DATA_TEMPR16[48] ), .B(\R_DATA_TEMPR17[48] ), 
        .C(\R_DATA_TEMPR18[48] ), .D(\R_DATA_TEMPR19[48] ), .Y(
        OR4_587_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%27%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C1 (
        .A_DOUT({\R_DATA_TEMPR27[79] , \R_DATA_TEMPR27[78] , 
        \R_DATA_TEMPR27[77] , \R_DATA_TEMPR27[76] , 
        \R_DATA_TEMPR27[75] , \R_DATA_TEMPR27[74] , 
        \R_DATA_TEMPR27[73] , \R_DATA_TEMPR27[72] , 
        \R_DATA_TEMPR27[71] , \R_DATA_TEMPR27[70] , 
        \R_DATA_TEMPR27[69] , \R_DATA_TEMPR27[68] , 
        \R_DATA_TEMPR27[67] , \R_DATA_TEMPR27[66] , 
        \R_DATA_TEMPR27[65] , \R_DATA_TEMPR27[64] , 
        \R_DATA_TEMPR27[63] , \R_DATA_TEMPR27[62] , 
        \R_DATA_TEMPR27[61] , \R_DATA_TEMPR27[60] }), .B_DOUT({
        \R_DATA_TEMPR27[59] , \R_DATA_TEMPR27[58] , 
        \R_DATA_TEMPR27[57] , \R_DATA_TEMPR27[56] , 
        \R_DATA_TEMPR27[55] , \R_DATA_TEMPR27[54] , 
        \R_DATA_TEMPR27[53] , \R_DATA_TEMPR27[52] , 
        \R_DATA_TEMPR27[51] , \R_DATA_TEMPR27[50] , 
        \R_DATA_TEMPR27[49] , \R_DATA_TEMPR27[48] , 
        \R_DATA_TEMPR27[47] , \R_DATA_TEMPR27[46] , 
        \R_DATA_TEMPR27[45] , \R_DATA_TEMPR27[44] , 
        \R_DATA_TEMPR27[43] , \R_DATA_TEMPR27[42] , 
        \R_DATA_TEMPR27[41] , \R_DATA_TEMPR27[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[27][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[6] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_545 (.A(\R_DATA_TEMPR8[47] ), .B(\R_DATA_TEMPR9[47] ), .C(
        \R_DATA_TEMPR10[47] ), .D(\R_DATA_TEMPR11[47] ), .Y(OR4_545_Y));
    OR4 OR4_233 (.A(OR4_390_Y), .B(OR2_20_Y), .C(\R_DATA_TEMPR22[66] ), 
        .D(\R_DATA_TEMPR23[66] ), .Y(OR4_233_Y));
    OR4 \OR4_R_DATA[41]  (.A(OR4_378_Y), .B(OR4_341_Y), .C(OR4_352_Y), 
        .D(OR4_120_Y), .Y(R_DATA[41]));
    OR4 OR4_562 (.A(OR4_506_Y), .B(OR4_351_Y), .C(OR4_513_Y), .D(
        OR4_109_Y), .Y(OR4_562_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%3%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0 (
        .A_DOUT({\R_DATA_TEMPR3[39] , \R_DATA_TEMPR3[38] , 
        \R_DATA_TEMPR3[37] , \R_DATA_TEMPR3[36] , \R_DATA_TEMPR3[35] , 
        \R_DATA_TEMPR3[34] , \R_DATA_TEMPR3[33] , \R_DATA_TEMPR3[32] , 
        \R_DATA_TEMPR3[31] , \R_DATA_TEMPR3[30] , \R_DATA_TEMPR3[29] , 
        \R_DATA_TEMPR3[28] , \R_DATA_TEMPR3[27] , \R_DATA_TEMPR3[26] , 
        \R_DATA_TEMPR3[25] , \R_DATA_TEMPR3[24] , \R_DATA_TEMPR3[23] , 
        \R_DATA_TEMPR3[22] , \R_DATA_TEMPR3[21] , \R_DATA_TEMPR3[20] })
        , .B_DOUT({\R_DATA_TEMPR3[19] , \R_DATA_TEMPR3[18] , 
        \R_DATA_TEMPR3[17] , \R_DATA_TEMPR3[16] , \R_DATA_TEMPR3[15] , 
        \R_DATA_TEMPR3[14] , \R_DATA_TEMPR3[13] , \R_DATA_TEMPR3[12] , 
        \R_DATA_TEMPR3[11] , \R_DATA_TEMPR3[10] , \R_DATA_TEMPR3[9] , 
        \R_DATA_TEMPR3[8] , \R_DATA_TEMPR3[7] , \R_DATA_TEMPR3[6] , 
        \R_DATA_TEMPR3[5] , \R_DATA_TEMPR3[4] , \R_DATA_TEMPR3[3] , 
        \R_DATA_TEMPR3[2] , \R_DATA_TEMPR3[1] , \R_DATA_TEMPR3[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[3][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_689 (.A(OR4_467_Y), .B(OR4_313_Y), .C(OR4_212_Y), .D(
        OR4_244_Y), .Y(OR4_689_Y));
    OR4 OR4_643 (.A(\R_DATA_TEMPR4[51] ), .B(\R_DATA_TEMPR5[51] ), .C(
        \R_DATA_TEMPR6[51] ), .D(\R_DATA_TEMPR7[51] ), .Y(OR4_643_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%12%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0 (
        .A_DOUT({\R_DATA_TEMPR12[39] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR12[37] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR12[35] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR12[33] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR12[31] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR12[29] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR12[27] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR12[25] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR12[23] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR12[21] , \R_DATA_TEMPR12[20] }), .B_DOUT({
        \R_DATA_TEMPR12[19] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR12[17] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR12[15] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR12[13] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR12[11] , \R_DATA_TEMPR12[10] , 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR12[8] , \R_DATA_TEMPR12[7] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR12[5] , \R_DATA_TEMPR12[4] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR12[2] , \R_DATA_TEMPR12[1] , 
        \R_DATA_TEMPR12[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_286 (.A(OR4_606_Y), .B(OR2_7_Y), .C(\R_DATA_TEMPR22[69] ), 
        .D(\R_DATA_TEMPR23[69] ), .Y(OR4_286_Y));
    OR4 OR4_78 (.A(\R_DATA_TEMPR0[4] ), .B(\R_DATA_TEMPR1[4] ), .C(
        \R_DATA_TEMPR2[4] ), .D(\R_DATA_TEMPR3[4] ), .Y(OR4_78_Y));
    OR4 \OR4_R_DATA[40]  (.A(OR4_256_Y), .B(OR4_403_Y), .C(OR4_10_Y), 
        .D(OR4_454_Y), .Y(R_DATA[40]));
    OR4 \OR4_R_DATA[8]  (.A(OR4_362_Y), .B(OR4_441_Y), .C(OR4_275_Y), 
        .D(OR4_542_Y), .Y(R_DATA[8]));
    OR4 OR4_564 (.A(OR4_190_Y), .B(OR2_1_Y), .C(\R_DATA_TEMPR22[78] ), 
        .D(\R_DATA_TEMPR23[78] ), .Y(OR4_564_Y));
    OR4 OR4_154 (.A(OR4_223_Y), .B(OR4_614_Y), .C(OR4_167_Y), .D(
        OR4_512_Y), .Y(OR4_154_Y));
    OR4 \OR4_R_DATA[61]  (.A(OR4_230_Y), .B(OR4_193_Y), .C(OR4_210_Y), 
        .D(OR4_697_Y), .Y(R_DATA[61]));
    OR4 OR4_684 (.A(\R_DATA_TEMPR0[16] ), .B(\R_DATA_TEMPR1[16] ), .C(
        \R_DATA_TEMPR2[16] ), .D(\R_DATA_TEMPR3[16] ), .Y(OR4_684_Y));
    OR2 OR2_21 (.A(\R_DATA_TEMPR20[3] ), .B(\R_DATA_TEMPR21[3] ), .Y(
        OR2_21_Y));
    OR4 OR4_638 (.A(\R_DATA_TEMPR0[38] ), .B(\R_DATA_TEMPR1[38] ), .C(
        \R_DATA_TEMPR2[38] ), .D(\R_DATA_TEMPR3[38] ), .Y(OR4_638_Y));
    OR4 OR4_22 (.A(\R_DATA_TEMPR8[41] ), .B(\R_DATA_TEMPR9[41] ), .C(
        \R_DATA_TEMPR10[41] ), .D(\R_DATA_TEMPR11[41] ), .Y(OR4_22_Y));
    OR2 OR2_73 (.A(\R_DATA_TEMPR20[75] ), .B(\R_DATA_TEMPR21[75] ), .Y(
        OR2_73_Y));
    OR4 \OR4_R_DATA[46]  (.A(OR4_713_Y), .B(OR4_381_Y), .C(OR4_510_Y), 
        .D(OR4_548_Y), .Y(R_DATA[46]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%29%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0 (
        .A_DOUT({\R_DATA_TEMPR29[39] , \R_DATA_TEMPR29[38] , 
        \R_DATA_TEMPR29[37] , \R_DATA_TEMPR29[36] , 
        \R_DATA_TEMPR29[35] , \R_DATA_TEMPR29[34] , 
        \R_DATA_TEMPR29[33] , \R_DATA_TEMPR29[32] , 
        \R_DATA_TEMPR29[31] , \R_DATA_TEMPR29[30] , 
        \R_DATA_TEMPR29[29] , \R_DATA_TEMPR29[28] , 
        \R_DATA_TEMPR29[27] , \R_DATA_TEMPR29[26] , 
        \R_DATA_TEMPR29[25] , \R_DATA_TEMPR29[24] , 
        \R_DATA_TEMPR29[23] , \R_DATA_TEMPR29[22] , 
        \R_DATA_TEMPR29[21] , \R_DATA_TEMPR29[20] }), .B_DOUT({
        \R_DATA_TEMPR29[19] , \R_DATA_TEMPR29[18] , 
        \R_DATA_TEMPR29[17] , \R_DATA_TEMPR29[16] , 
        \R_DATA_TEMPR29[15] , \R_DATA_TEMPR29[14] , 
        \R_DATA_TEMPR29[13] , \R_DATA_TEMPR29[12] , 
        \R_DATA_TEMPR29[11] , \R_DATA_TEMPR29[10] , 
        \R_DATA_TEMPR29[9] , \R_DATA_TEMPR29[8] , \R_DATA_TEMPR29[7] , 
        \R_DATA_TEMPR29[6] , \R_DATA_TEMPR29[5] , \R_DATA_TEMPR29[4] , 
        \R_DATA_TEMPR29[3] , \R_DATA_TEMPR29[2] , \R_DATA_TEMPR29[1] , 
        \R_DATA_TEMPR29[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_143 (.A(\R_DATA_TEMPR12[8] ), .B(\R_DATA_TEMPR13[8] ), .C(
        \R_DATA_TEMPR14[8] ), .D(\R_DATA_TEMPR15[8] ), .Y(OR4_143_Y));
    OR4 OR4_632 (.A(\R_DATA_TEMPR24[50] ), .B(\R_DATA_TEMPR25[50] ), 
        .C(\R_DATA_TEMPR26[50] ), .D(\R_DATA_TEMPR27[50] ), .Y(
        OR4_632_Y));
    OR4 OR4_213 (.A(\R_DATA_TEMPR24[73] ), .B(\R_DATA_TEMPR25[73] ), 
        .C(\R_DATA_TEMPR26[73] ), .D(\R_DATA_TEMPR27[73] ), .Y(
        OR4_213_Y));
    OR4 OR4_201 (.A(\R_DATA_TEMPR4[43] ), .B(\R_DATA_TEMPR5[43] ), .C(
        \R_DATA_TEMPR6[43] ), .D(\R_DATA_TEMPR7[43] ), .Y(OR4_201_Y));
    OR4 OR4_361 (.A(\R_DATA_TEMPR28[18] ), .B(\R_DATA_TEMPR29[18] ), 
        .C(\R_DATA_TEMPR30[18] ), .D(\R_DATA_TEMPR31[18] ), .Y(
        OR4_361_Y));
    OR4 \OR4_R_DATA[74]  (.A(OR4_660_Y), .B(OR4_402_Y), .C(OR4_39_Y), 
        .D(OR4_348_Y), .Y(R_DATA[74]));
    OR4 \OR4_R_DATA[60]  (.A(OR4_81_Y), .B(OR4_263_Y), .C(OR4_578_Y), 
        .D(OR4_299_Y), .Y(R_DATA[60]));
    OR2 OR2_13 (.A(\R_DATA_TEMPR20[5] ), .B(\R_DATA_TEMPR21[5] ), .Y(
        OR2_13_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%21%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0 (
        .A_DOUT({\R_DATA_TEMPR21[39] , \R_DATA_TEMPR21[38] , 
        \R_DATA_TEMPR21[37] , \R_DATA_TEMPR21[36] , 
        \R_DATA_TEMPR21[35] , \R_DATA_TEMPR21[34] , 
        \R_DATA_TEMPR21[33] , \R_DATA_TEMPR21[32] , 
        \R_DATA_TEMPR21[31] , \R_DATA_TEMPR21[30] , 
        \R_DATA_TEMPR21[29] , \R_DATA_TEMPR21[28] , 
        \R_DATA_TEMPR21[27] , \R_DATA_TEMPR21[26] , 
        \R_DATA_TEMPR21[25] , \R_DATA_TEMPR21[24] , 
        \R_DATA_TEMPR21[23] , \R_DATA_TEMPR21[22] , 
        \R_DATA_TEMPR21[21] , \R_DATA_TEMPR21[20] }), .B_DOUT({
        \R_DATA_TEMPR21[19] , \R_DATA_TEMPR21[18] , 
        \R_DATA_TEMPR21[17] , \R_DATA_TEMPR21[16] , 
        \R_DATA_TEMPR21[15] , \R_DATA_TEMPR21[14] , 
        \R_DATA_TEMPR21[13] , \R_DATA_TEMPR21[12] , 
        \R_DATA_TEMPR21[11] , \R_DATA_TEMPR21[10] , 
        \R_DATA_TEMPR21[9] , \R_DATA_TEMPR21[8] , \R_DATA_TEMPR21[7] , 
        \R_DATA_TEMPR21[6] , \R_DATA_TEMPR21[5] , \R_DATA_TEMPR21[4] , 
        \R_DATA_TEMPR21[3] , \R_DATA_TEMPR21[2] , \R_DATA_TEMPR21[1] , 
        \R_DATA_TEMPR21[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_6 (.A(OR4_182_Y), .B(OR2_67_Y), .C(\R_DATA_TEMPR22[16] ), 
        .D(\R_DATA_TEMPR23[16] ), .Y(OR4_6_Y));
    OR4 OR4_271 (.A(\R_DATA_TEMPR4[45] ), .B(\R_DATA_TEMPR5[45] ), .C(
        \R_DATA_TEMPR6[45] ), .D(\R_DATA_TEMPR7[45] ), .Y(OR4_271_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%24%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C1 (
        .A_DOUT({\R_DATA_TEMPR24[79] , \R_DATA_TEMPR24[78] , 
        \R_DATA_TEMPR24[77] , \R_DATA_TEMPR24[76] , 
        \R_DATA_TEMPR24[75] , \R_DATA_TEMPR24[74] , 
        \R_DATA_TEMPR24[73] , \R_DATA_TEMPR24[72] , 
        \R_DATA_TEMPR24[71] , \R_DATA_TEMPR24[70] , 
        \R_DATA_TEMPR24[69] , \R_DATA_TEMPR24[68] , 
        \R_DATA_TEMPR24[67] , \R_DATA_TEMPR24[66] , 
        \R_DATA_TEMPR24[65] , \R_DATA_TEMPR24[64] , 
        \R_DATA_TEMPR24[63] , \R_DATA_TEMPR24[62] , 
        \R_DATA_TEMPR24[61] , \R_DATA_TEMPR24[60] }), .B_DOUT({
        \R_DATA_TEMPR24[59] , \R_DATA_TEMPR24[58] , 
        \R_DATA_TEMPR24[57] , \R_DATA_TEMPR24[56] , 
        \R_DATA_TEMPR24[55] , \R_DATA_TEMPR24[54] , 
        \R_DATA_TEMPR24[53] , \R_DATA_TEMPR24[52] , 
        \R_DATA_TEMPR24[51] , \R_DATA_TEMPR24[50] , 
        \R_DATA_TEMPR24[49] , \R_DATA_TEMPR24[48] , 
        \R_DATA_TEMPR24[47] , \R_DATA_TEMPR24[46] , 
        \R_DATA_TEMPR24[45] , \R_DATA_TEMPR24[44] , 
        \R_DATA_TEMPR24[43] , \R_DATA_TEMPR24[42] , 
        \R_DATA_TEMPR24[41] , \R_DATA_TEMPR24[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[24][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_460 (.A(\R_DATA_TEMPR12[63] ), .B(\R_DATA_TEMPR13[63] ), 
        .C(\R_DATA_TEMPR14[63] ), .D(\R_DATA_TEMPR15[63] ), .Y(
        OR4_460_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%28%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0 (
        .A_DOUT({\R_DATA_TEMPR28[39] , \R_DATA_TEMPR28[38] , 
        \R_DATA_TEMPR28[37] , \R_DATA_TEMPR28[36] , 
        \R_DATA_TEMPR28[35] , \R_DATA_TEMPR28[34] , 
        \R_DATA_TEMPR28[33] , \R_DATA_TEMPR28[32] , 
        \R_DATA_TEMPR28[31] , \R_DATA_TEMPR28[30] , 
        \R_DATA_TEMPR28[29] , \R_DATA_TEMPR28[28] , 
        \R_DATA_TEMPR28[27] , \R_DATA_TEMPR28[26] , 
        \R_DATA_TEMPR28[25] , \R_DATA_TEMPR28[24] , 
        \R_DATA_TEMPR28[23] , \R_DATA_TEMPR28[22] , 
        \R_DATA_TEMPR28[21] , \R_DATA_TEMPR28[20] }), .B_DOUT({
        \R_DATA_TEMPR28[19] , \R_DATA_TEMPR28[18] , 
        \R_DATA_TEMPR28[17] , \R_DATA_TEMPR28[16] , 
        \R_DATA_TEMPR28[15] , \R_DATA_TEMPR28[14] , 
        \R_DATA_TEMPR28[13] , \R_DATA_TEMPR28[12] , 
        \R_DATA_TEMPR28[11] , \R_DATA_TEMPR28[10] , 
        \R_DATA_TEMPR28[9] , \R_DATA_TEMPR28[8] , \R_DATA_TEMPR28[7] , 
        \R_DATA_TEMPR28[6] , \R_DATA_TEMPR28[5] , \R_DATA_TEMPR28[4] , 
        \R_DATA_TEMPR28[3] , \R_DATA_TEMPR28[2] , \R_DATA_TEMPR28[1] , 
        \R_DATA_TEMPR28[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_502 (.A(OR4_209_Y), .B(OR2_4_Y), .C(\R_DATA_TEMPR22[12] ), 
        .D(\R_DATA_TEMPR23[12] ), .Y(OR4_502_Y));
    OR4 \OR4_R_DATA[66]  (.A(OR4_558_Y), .B(OR4_233_Y), .C(OR4_350_Y), 
        .D(OR4_388_Y), .Y(R_DATA[66]));
    OR4 OR4_556 (.A(OR4_78_Y), .B(OR4_225_Y), .C(OR4_86_Y), .D(
        OR4_463_Y), .Y(OR4_556_Y));
    OR4 OR4_495 (.A(OR4_626_Y), .B(OR4_322_Y), .C(OR4_486_Y), .D(
        OR4_108_Y), .Y(OR4_495_Y));
    OR4 OR4_572 (.A(\R_DATA_TEMPR0[14] ), .B(\R_DATA_TEMPR1[14] ), .C(
        \R_DATA_TEMPR2[14] ), .D(\R_DATA_TEMPR3[14] ), .Y(OR4_572_Y));
    OR2 OR2_54 (.A(\R_DATA_TEMPR20[59] ), .B(\R_DATA_TEMPR21[59] ), .Y(
        OR2_54_Y));
    OR4 OR4_618 (.A(\R_DATA_TEMPR24[62] ), .B(\R_DATA_TEMPR25[62] ), 
        .C(\R_DATA_TEMPR26[62] ), .D(\R_DATA_TEMPR27[62] ), .Y(
        OR4_618_Y));
    OR2 OR2_71 (.A(\R_DATA_TEMPR20[27] ), .B(\R_DATA_TEMPR21[27] ), .Y(
        OR2_71_Y));
    OR4 \OR4_R_DATA[17]  (.A(OR4_154_Y), .B(OR4_501_Y), .C(OR4_682_Y), 
        .D(OR4_29_Y), .Y(R_DATA[17]));
    OR4 OR4_142 (.A(\R_DATA_TEMPR24[31] ), .B(\R_DATA_TEMPR25[31] ), 
        .C(\R_DATA_TEMPR26[31] ), .D(\R_DATA_TEMPR27[31] ), .Y(
        OR4_142_Y));
    OR4 OR4_612 (.A(\R_DATA_TEMPR4[15] ), .B(\R_DATA_TEMPR5[15] ), .C(
        \R_DATA_TEMPR6[15] ), .D(\R_DATA_TEMPR7[15] ), .Y(OR4_612_Y));
    OR4 OR4_504 (.A(OR4_121_Y), .B(OR4_644_Y), .C(OR4_676_Y), .D(
        OR4_73_Y), .Y(OR4_504_Y));
    OR4 OR4_574 (.A(\R_DATA_TEMPR8[48] ), .B(\R_DATA_TEMPR9[48] ), .C(
        \R_DATA_TEMPR10[48] ), .D(\R_DATA_TEMPR11[48] ), .Y(OR4_574_Y));
    OR2 OR2_11 (.A(\R_DATA_TEMPR20[50] ), .B(\R_DATA_TEMPR21[50] ), .Y(
        OR2_11_Y));
    OR4 OR4_494 (.A(\R_DATA_TEMPR28[35] ), .B(\R_DATA_TEMPR29[35] ), 
        .C(\R_DATA_TEMPR30[35] ), .D(\R_DATA_TEMPR31[35] ), .Y(
        OR4_494_Y));
    OR4 OR4_558 (.A(OR4_188_Y), .B(OR4_687_Y), .C(OR4_1_Y), .D(
        OR4_124_Y), .Y(OR4_558_Y));
    OR4 OR4_55 (.A(\R_DATA_TEMPR12[57] ), .B(\R_DATA_TEMPR13[57] ), .C(
        \R_DATA_TEMPR14[57] ), .D(\R_DATA_TEMPR15[57] ), .Y(OR4_55_Y));
    OR4 OR4_369 (.A(OR4_426_Y), .B(OR4_95_Y), .C(OR4_385_Y), .D(
        OR4_5_Y), .Y(OR4_369_Y));
    OR4 OR4_301 (.A(\R_DATA_TEMPR24[20] ), .B(\R_DATA_TEMPR25[20] ), 
        .C(\R_DATA_TEMPR26[20] ), .D(\R_DATA_TEMPR27[20] ), .Y(
        OR4_301_Y));
    OR4 OR4_396 (.A(\R_DATA_TEMPR12[38] ), .B(\R_DATA_TEMPR13[38] ), 
        .C(\R_DATA_TEMPR14[38] ), .D(\R_DATA_TEMPR15[38] ), .Y(
        OR4_396_Y));
    OR4 OR4_249 (.A(OR4_12_Y), .B(OR4_588_Y), .C(OR4_465_Y), .D(
        OR4_500_Y), .Y(OR4_249_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%1%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0 (
        .A_DOUT({\R_DATA_TEMPR1[39] , \R_DATA_TEMPR1[38] , 
        \R_DATA_TEMPR1[37] , \R_DATA_TEMPR1[36] , \R_DATA_TEMPR1[35] , 
        \R_DATA_TEMPR1[34] , \R_DATA_TEMPR1[33] , \R_DATA_TEMPR1[32] , 
        \R_DATA_TEMPR1[31] , \R_DATA_TEMPR1[30] , \R_DATA_TEMPR1[29] , 
        \R_DATA_TEMPR1[28] , \R_DATA_TEMPR1[27] , \R_DATA_TEMPR1[26] , 
        \R_DATA_TEMPR1[25] , \R_DATA_TEMPR1[24] , \R_DATA_TEMPR1[23] , 
        \R_DATA_TEMPR1[22] , \R_DATA_TEMPR1[21] , \R_DATA_TEMPR1[20] })
        , .B_DOUT({\R_DATA_TEMPR1[19] , \R_DATA_TEMPR1[18] , 
        \R_DATA_TEMPR1[17] , \R_DATA_TEMPR1[16] , \R_DATA_TEMPR1[15] , 
        \R_DATA_TEMPR1[14] , \R_DATA_TEMPR1[13] , \R_DATA_TEMPR1[12] , 
        \R_DATA_TEMPR1[11] , \R_DATA_TEMPR1[10] , \R_DATA_TEMPR1[9] , 
        \R_DATA_TEMPR1[8] , \R_DATA_TEMPR1[7] , \R_DATA_TEMPR1[6] , 
        \R_DATA_TEMPR1[5] , \R_DATA_TEMPR1[4] , \R_DATA_TEMPR1[3] , 
        \R_DATA_TEMPR1[2] , \R_DATA_TEMPR1[1] , \R_DATA_TEMPR1[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[1][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_371 (.A(\R_DATA_TEMPR28[3] ), .B(\R_DATA_TEMPR29[3] ), .C(
        \R_DATA_TEMPR30[3] ), .D(\R_DATA_TEMPR31[3] ), .Y(OR4_371_Y));
    OR4 OR4_425 (.A(\R_DATA_TEMPR24[38] ), .B(\R_DATA_TEMPR25[38] ), 
        .C(\R_DATA_TEMPR26[38] ), .D(\R_DATA_TEMPR27[38] ), .Y(
        OR4_425_Y));
    OR4 OR4_400 (.A(\R_DATA_TEMPR28[47] ), .B(\R_DATA_TEMPR29[47] ), 
        .C(\R_DATA_TEMPR30[47] ), .D(\R_DATA_TEMPR31[47] ), .Y(
        OR4_400_Y));
    OR4 OR4_636 (.A(OR4_204_Y), .B(OR4_612_Y), .C(OR4_646_Y), .D(
        OR4_284_Y), .Y(OR4_636_Y));
    OR4 \OR4_R_DATA[38]  (.A(OR4_125_Y), .B(OR4_38_Y), .C(OR4_425_Y), 
        .D(OR4_531_Y), .Y(R_DATA[38]));
    OR4 OR4_456 (.A(\R_DATA_TEMPR0[55] ), .B(\R_DATA_TEMPR1[55] ), .C(
        \R_DATA_TEMPR2[55] ), .D(\R_DATA_TEMPR3[55] ), .Y(OR4_456_Y));
    OR4 OR4_470 (.A(\R_DATA_TEMPR28[53] ), .B(\R_DATA_TEMPR29[53] ), 
        .C(\R_DATA_TEMPR30[53] ), .D(\R_DATA_TEMPR31[53] ), .Y(
        OR4_470_Y));
    OR4 \OR4_R_DATA[47]  (.A(OR4_530_Y), .B(OR4_153_Y), .C(OR4_329_Y), 
        .D(OR4_400_Y), .Y(R_DATA[47]));
    OR4 OR4_352 (.A(\R_DATA_TEMPR24[41] ), .B(\R_DATA_TEMPR25[41] ), 
        .C(\R_DATA_TEMPR26[41] ), .D(\R_DATA_TEMPR27[41] ), .Y(
        OR4_352_Y));
    OR4 OR4_15 (.A(\R_DATA_TEMPR0[69] ), .B(\R_DATA_TEMPR1[69] ), .C(
        \R_DATA_TEMPR2[69] ), .D(\R_DATA_TEMPR3[69] ), .Y(OR4_15_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[3]  (.A(CFG2_0_Y), .B(
        W_ADDR[13]), .C(W_EN), .Y(\BLKX2[3] ));
    OR4 OR4_424 (.A(\R_DATA_TEMPR16[68] ), .B(\R_DATA_TEMPR17[68] ), 
        .C(\R_DATA_TEMPR18[68] ), .D(\R_DATA_TEMPR19[68] ), .Y(
        OR4_424_Y));
    OR4 OR4_281 (.A(\R_DATA_TEMPR16[44] ), .B(\R_DATA_TEMPR17[44] ), 
        .C(\R_DATA_TEMPR18[44] ), .D(\R_DATA_TEMPR19[44] ), .Y(
        OR4_281_Y));
    OR4 OR4_194 (.A(\R_DATA_TEMPR24[45] ), .B(\R_DATA_TEMPR25[45] ), 
        .C(\R_DATA_TEMPR26[45] ), .D(\R_DATA_TEMPR27[45] ), .Y(
        OR4_194_Y));
    OR4 \OR4_R_DATA[67]  (.A(OR4_369_Y), .B(OR4_715_Y), .C(OR4_186_Y), 
        .D(OR4_257_Y), .Y(R_DATA[67]));
    OR4 OR4_326 (.A(\R_DATA_TEMPR28[78] ), .B(\R_DATA_TEMPR29[78] ), 
        .C(\R_DATA_TEMPR30[78] ), .D(\R_DATA_TEMPR31[78] ), .Y(
        OR4_326_Y));
    OR4 OR4_563 (.A(\R_DATA_TEMPR16[37] ), .B(\R_DATA_TEMPR17[37] ), 
        .C(\R_DATA_TEMPR18[37] ), .D(\R_DATA_TEMPR19[37] ), .Y(
        OR4_563_Y));
    OR4 OR4_93 (.A(\R_DATA_TEMPR12[64] ), .B(\R_DATA_TEMPR13[64] ), .C(
        \R_DATA_TEMPR14[64] ), .D(\R_DATA_TEMPR15[64] ), .Y(OR4_93_Y));
    OR4 OR4_616 (.A(\R_DATA_TEMPR16[67] ), .B(\R_DATA_TEMPR17[67] ), 
        .C(\R_DATA_TEMPR18[67] ), .D(\R_DATA_TEMPR19[67] ), .Y(
        OR4_616_Y));
    OR4 OR4_309 (.A(OR4_659_Y), .B(OR4_438_Y), .C(OR4_487_Y), .D(
        OR4_613_Y), .Y(OR4_309_Y));
    OR4 OR4_582 (.A(\R_DATA_TEMPR8[25] ), .B(\R_DATA_TEMPR9[25] ), .C(
        \R_DATA_TEMPR10[25] ), .D(\R_DATA_TEMPR11[25] ), .Y(OR4_582_Y));
    OR4 OR4_24 (.A(\R_DATA_TEMPR24[19] ), .B(\R_DATA_TEMPR25[19] ), .C(
        \R_DATA_TEMPR26[19] ), .D(\R_DATA_TEMPR27[19] ), .Y(OR4_24_Y));
    OR4 OR4_8 (.A(\R_DATA_TEMPR4[42] ), .B(\R_DATA_TEMPR5[42] ), .C(
        \R_DATA_TEMPR6[42] ), .D(\R_DATA_TEMPR7[42] ), .Y(OR4_8_Y));
    OR4 OR4_379 (.A(\R_DATA_TEMPR0[37] ), .B(\R_DATA_TEMPR1[37] ), .C(
        \R_DATA_TEMPR2[37] ), .D(\R_DATA_TEMPR3[37] ), .Y(OR4_379_Y));
    OR4 OR4_250 (.A(OR4_442_Y), .B(OR2_31_Y), .C(\R_DATA_TEMPR22[51] ), 
        .D(\R_DATA_TEMPR23[51] ), .Y(OR4_250_Y));
    OR4 OR4_557 (.A(\R_DATA_TEMPR12[55] ), .B(\R_DATA_TEMPR13[55] ), 
        .C(\R_DATA_TEMPR14[55] ), .D(\R_DATA_TEMPR15[55] ), .Y(
        OR4_557_Y));
    OR2 OR2_4 (.A(\R_DATA_TEMPR20[12] ), .B(\R_DATA_TEMPR21[12] ), .Y(
        OR2_4_Y));
    OR4 OR4_334 (.A(\R_DATA_TEMPR0[46] ), .B(\R_DATA_TEMPR1[46] ), .C(
        \R_DATA_TEMPR2[46] ), .D(\R_DATA_TEMPR3[46] ), .Y(OR4_334_Y));
    OR4 \OR4_R_DATA[71]  (.A(OR4_700_Y), .B(OR4_664_Y), .C(OR4_674_Y), 
        .D(OR4_447_Y), .Y(R_DATA[71]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%18%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C1 (
        .A_DOUT({\R_DATA_TEMPR18[79] , \R_DATA_TEMPR18[78] , 
        \R_DATA_TEMPR18[77] , \R_DATA_TEMPR18[76] , 
        \R_DATA_TEMPR18[75] , \R_DATA_TEMPR18[74] , 
        \R_DATA_TEMPR18[73] , \R_DATA_TEMPR18[72] , 
        \R_DATA_TEMPR18[71] , \R_DATA_TEMPR18[70] , 
        \R_DATA_TEMPR18[69] , \R_DATA_TEMPR18[68] , 
        \R_DATA_TEMPR18[67] , \R_DATA_TEMPR18[66] , 
        \R_DATA_TEMPR18[65] , \R_DATA_TEMPR18[64] , 
        \R_DATA_TEMPR18[63] , \R_DATA_TEMPR18[62] , 
        \R_DATA_TEMPR18[61] , \R_DATA_TEMPR18[60] }), .B_DOUT({
        \R_DATA_TEMPR18[59] , \R_DATA_TEMPR18[58] , 
        \R_DATA_TEMPR18[57] , \R_DATA_TEMPR18[56] , 
        \R_DATA_TEMPR18[55] , \R_DATA_TEMPR18[54] , 
        \R_DATA_TEMPR18[53] , \R_DATA_TEMPR18[52] , 
        \R_DATA_TEMPR18[51] , \R_DATA_TEMPR18[50] , 
        \R_DATA_TEMPR18[49] , \R_DATA_TEMPR18[48] , 
        \R_DATA_TEMPR18[47] , \R_DATA_TEMPR18[46] , 
        \R_DATA_TEMPR18[45] , \R_DATA_TEMPR18[44] , 
        \R_DATA_TEMPR18[43] , \R_DATA_TEMPR18[42] , 
        \R_DATA_TEMPR18[41] , \R_DATA_TEMPR18[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[18][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[4] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_131 (.A(OR4_72_Y), .B(OR4_651_Y), .C(OR4_79_Y), .D(
        OR4_414_Y), .Y(OR4_131_Y));
    OR4 OR4_584 (.A(\R_DATA_TEMPR4[77] ), .B(\R_DATA_TEMPR5[77] ), .C(
        \R_DATA_TEMPR6[77] ), .D(\R_DATA_TEMPR7[77] ), .Y(OR4_584_Y));
    OR4 OR4_659 (.A(\R_DATA_TEMPR0[76] ), .B(\R_DATA_TEMPR1[76] ), .C(
        \R_DATA_TEMPR2[76] ), .D(\R_DATA_TEMPR3[76] ), .Y(OR4_659_Y));
    OR4 OR4_596 (.A(\R_DATA_TEMPR0[22] ), .B(\R_DATA_TEMPR1[22] ), .C(
        \R_DATA_TEMPR2[22] ), .D(\R_DATA_TEMPR3[22] ), .Y(OR4_596_Y));
    OR4 \OR4_R_DATA[39]  (.A(OR4_393_Y), .B(OR4_252_Y), .C(OR4_202_Y), 
        .D(OR4_58_Y), .Y(R_DATA[39]));
    OR4 OR4_256 (.A(OR4_199_Y), .B(OR4_35_Y), .C(OR4_207_Y), .D(
        OR4_523_Y), .Y(OR4_256_Y));
    OR2 OR2_0 (.A(\R_DATA_TEMPR20[74] ), .B(\R_DATA_TEMPR21[74] ), .Y(
        OR2_0_Y));
    OR4 OR4_75 (.A(\R_DATA_TEMPR4[53] ), .B(\R_DATA_TEMPR5[53] ), .C(
        \R_DATA_TEMPR6[53] ), .D(\R_DATA_TEMPR7[53] ), .Y(OR4_75_Y));
    OR2 OR2_6 (.A(\R_DATA_TEMPR20[33] ), .B(\R_DATA_TEMPR21[33] ), .Y(
        OR2_6_Y));
    OR4 OR4_431 (.A(\R_DATA_TEMPR28[56] ), .B(\R_DATA_TEMPR29[56] ), 
        .C(\R_DATA_TEMPR30[56] ), .D(\R_DATA_TEMPR31[56] ), .Y(
        OR4_431_Y));
    OR4 \OR4_R_DATA[70]  (.A(OR4_562_Y), .B(OR4_3_Y), .C(OR4_323_Y), 
        .D(OR4_54_Y), .Y(R_DATA[70]));
    OR4 OR4_91 (.A(\R_DATA_TEMPR0[32] ), .B(\R_DATA_TEMPR1[32] ), .C(
        \R_DATA_TEMPR2[32] ), .D(\R_DATA_TEMPR3[32] ), .Y(OR4_91_Y));
    OR4 OR4_124 (.A(\R_DATA_TEMPR12[66] ), .B(\R_DATA_TEMPR13[66] ), 
        .C(\R_DATA_TEMPR14[66] ), .D(\R_DATA_TEMPR15[66] ), .Y(
        OR4_124_Y));
    OR4 OR4_438 (.A(\R_DATA_TEMPR4[76] ), .B(\R_DATA_TEMPR5[76] ), .C(
        \R_DATA_TEMPR6[76] ), .D(\R_DATA_TEMPR7[76] ), .Y(OR4_438_Y));
    OR4 OR4_709 (.A(\R_DATA_TEMPR4[33] ), .B(\R_DATA_TEMPR5[33] ), .C(
        \R_DATA_TEMPR6[33] ), .D(\R_DATA_TEMPR7[33] ), .Y(OR4_709_Y));
    OR4 OR4_381 (.A(OR4_553_Y), .B(OR2_59_Y), .C(\R_DATA_TEMPR22[46] ), 
        .D(\R_DATA_TEMPR23[46] ), .Y(OR4_381_Y));
    OR2 OR2_3 (.A(\R_DATA_TEMPR20[71] ), .B(\R_DATA_TEMPR21[71] ), .Y(
        OR2_3_Y));
    OR4 OR4_654 (.A(\R_DATA_TEMPR0[73] ), .B(\R_DATA_TEMPR1[73] ), .C(
        \R_DATA_TEMPR2[73] ), .D(\R_DATA_TEMPR3[73] ), .Y(OR4_654_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[5]  (.A(CFG2_2_Y), .B(
        W_ADDR[13]), .C(W_EN), .Y(\BLKX2[5] ));
    OR4 \OR4_R_DATA[76]  (.A(OR4_309_Y), .B(OR4_705_Y), .C(OR4_97_Y), 
        .D(OR4_141_Y), .Y(R_DATA[76]));
    OR4 OR4_480 (.A(\R_DATA_TEMPR24[1] ), .B(\R_DATA_TEMPR25[1] ), .C(
        \R_DATA_TEMPR26[1] ), .D(\R_DATA_TEMPR27[1] ), .Y(OR4_480_Y));
    OR4 OR4_503 (.A(\R_DATA_TEMPR12[65] ), .B(\R_DATA_TEMPR13[65] ), 
        .C(\R_DATA_TEMPR14[65] ), .D(\R_DATA_TEMPR15[65] ), .Y(
        OR4_503_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[7]  (.A(CFG2_0_Y), .B(
        W_ADDR[13]), .C(W_EN), .Y(\BLKX2[7] ));
    OR4 OR4_314 (.A(\R_DATA_TEMPR24[3] ), .B(\R_DATA_TEMPR25[3] ), .C(
        \R_DATA_TEMPR26[3] ), .D(\R_DATA_TEMPR27[3] ), .Y(OR4_314_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%20%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0 (
        .A_DOUT({\R_DATA_TEMPR20[39] , \R_DATA_TEMPR20[38] , 
        \R_DATA_TEMPR20[37] , \R_DATA_TEMPR20[36] , 
        \R_DATA_TEMPR20[35] , \R_DATA_TEMPR20[34] , 
        \R_DATA_TEMPR20[33] , \R_DATA_TEMPR20[32] , 
        \R_DATA_TEMPR20[31] , \R_DATA_TEMPR20[30] , 
        \R_DATA_TEMPR20[29] , \R_DATA_TEMPR20[28] , 
        \R_DATA_TEMPR20[27] , \R_DATA_TEMPR20[26] , 
        \R_DATA_TEMPR20[25] , \R_DATA_TEMPR20[24] , 
        \R_DATA_TEMPR20[23] , \R_DATA_TEMPR20[22] , 
        \R_DATA_TEMPR20[21] , \R_DATA_TEMPR20[20] }), .B_DOUT({
        \R_DATA_TEMPR20[19] , \R_DATA_TEMPR20[18] , 
        \R_DATA_TEMPR20[17] , \R_DATA_TEMPR20[16] , 
        \R_DATA_TEMPR20[15] , \R_DATA_TEMPR20[14] , 
        \R_DATA_TEMPR20[13] , \R_DATA_TEMPR20[12] , 
        \R_DATA_TEMPR20[11] , \R_DATA_TEMPR20[10] , 
        \R_DATA_TEMPR20[9] , \R_DATA_TEMPR20[8] , \R_DATA_TEMPR20[7] , 
        \R_DATA_TEMPR20[6] , \R_DATA_TEMPR20[5] , \R_DATA_TEMPR20[4] , 
        \R_DATA_TEMPR20[3] , \R_DATA_TEMPR20[2] , \R_DATA_TEMPR20[1] , 
        \R_DATA_TEMPR20[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_43 (.A(OR4_668_Y), .B(OR2_45_Y), .C(\R_DATA_TEMPR22[57] ), 
        .D(\R_DATA_TEMPR23[57] ), .Y(OR4_43_Y));
    OR4 OR4_573 (.A(\R_DATA_TEMPR0[0] ), .B(\R_DATA_TEMPR1[0] ), .C(
        \R_DATA_TEMPR2[0] ), .D(\R_DATA_TEMPR3[0] ), .Y(OR4_573_Y));
    OR4 OR4_539 (.A(\R_DATA_TEMPR0[10] ), .B(\R_DATA_TEMPR1[10] ), .C(
        \R_DATA_TEMPR2[10] ), .D(\R_DATA_TEMPR3[10] ), .Y(OR4_539_Y));
    INV \INVBLKX0[0]  (.A(W_ADDR[9]), .Y(\BLKX0[0] ));
    OR2 OR2_26 (.A(\R_DATA_TEMPR20[54] ), .B(\R_DATA_TEMPR21[54] ), .Y(
        OR2_26_Y));
    OR4 OR4_111 (.A(\R_DATA_TEMPR0[48] ), .B(\R_DATA_TEMPR1[48] ), .C(
        \R_DATA_TEMPR2[48] ), .D(\R_DATA_TEMPR3[48] ), .Y(OR4_111_Y));
    OR4 OR4_598 (.A(\R_DATA_TEMPR28[64] ), .B(\R_DATA_TEMPR29[64] ), 
        .C(\R_DATA_TEMPR30[64] ), .D(\R_DATA_TEMPR31[64] ), .Y(
        OR4_598_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%16%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C1 (
        .A_DOUT({\R_DATA_TEMPR16[79] , \R_DATA_TEMPR16[78] , 
        \R_DATA_TEMPR16[77] , \R_DATA_TEMPR16[76] , 
        \R_DATA_TEMPR16[75] , \R_DATA_TEMPR16[74] , 
        \R_DATA_TEMPR16[73] , \R_DATA_TEMPR16[72] , 
        \R_DATA_TEMPR16[71] , \R_DATA_TEMPR16[70] , 
        \R_DATA_TEMPR16[69] , \R_DATA_TEMPR16[68] , 
        \R_DATA_TEMPR16[67] , \R_DATA_TEMPR16[66] , 
        \R_DATA_TEMPR16[65] , \R_DATA_TEMPR16[64] , 
        \R_DATA_TEMPR16[63] , \R_DATA_TEMPR16[62] , 
        \R_DATA_TEMPR16[61] , \R_DATA_TEMPR16[60] }), .B_DOUT({
        \R_DATA_TEMPR16[59] , \R_DATA_TEMPR16[58] , 
        \R_DATA_TEMPR16[57] , \R_DATA_TEMPR16[56] , 
        \R_DATA_TEMPR16[55] , \R_DATA_TEMPR16[54] , 
        \R_DATA_TEMPR16[53] , \R_DATA_TEMPR16[52] , 
        \R_DATA_TEMPR16[51] , \R_DATA_TEMPR16[50] , 
        \R_DATA_TEMPR16[49] , \R_DATA_TEMPR16[48] , 
        \R_DATA_TEMPR16[47] , \R_DATA_TEMPR16[46] , 
        \R_DATA_TEMPR16[45] , \R_DATA_TEMPR16[44] , 
        \R_DATA_TEMPR16[43] , \R_DATA_TEMPR16[42] , 
        \R_DATA_TEMPR16[41] , \R_DATA_TEMPR16[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[16][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_59 (.A(\R_DATA_TEMPR0[64] ), .B(\R_DATA_TEMPR1[64] ), .C(
        \R_DATA_TEMPR2[64] ), .D(\R_DATA_TEMPR3[64] ), .Y(OR4_59_Y));
    OR4 OR4_530 (.A(OR4_591_Y), .B(OR4_273_Y), .C(OR4_545_Y), .D(
        OR4_162_Y), .Y(OR4_530_Y));
    OR4 OR4_263 (.A(OR4_355_Y), .B(OR2_50_Y), .C(\R_DATA_TEMPR22[60] ), 
        .D(\R_DATA_TEMPR23[60] ), .Y(OR4_263_Y));
    OR4 OR4_526 (.A(OR4_656_Y), .B(OR4_356_Y), .C(OR4_508_Y), .D(
        OR4_144_Y), .Y(OR4_526_Y));
    OR4 OR4_445 (.A(\R_DATA_TEMPR8[22] ), .B(\R_DATA_TEMPR9[22] ), .C(
        \R_DATA_TEMPR10[22] ), .D(\R_DATA_TEMPR11[22] ), .Y(OR4_445_Y));
    OR4 OR4_411 (.A(\R_DATA_TEMPR12[52] ), .B(\R_DATA_TEMPR13[52] ), 
        .C(\R_DATA_TEMPR14[52] ), .D(\R_DATA_TEMPR15[52] ), .Y(
        OR4_411_Y));
    OR4 OR4_496 (.A(\R_DATA_TEMPR16[43] ), .B(\R_DATA_TEMPR17[43] ), 
        .C(\R_DATA_TEMPR18[43] ), .D(\R_DATA_TEMPR19[43] ), .Y(
        OR4_496_Y));
    OR4 OR4_418 (.A(OR4_130_Y), .B(OR2_30_Y), .C(\R_DATA_TEMPR22[35] ), 
        .D(\R_DATA_TEMPR23[35] ), .Y(OR4_418_Y));
    OR4 \OR4_R_DATA[0]  (.A(OR4_599_Y), .B(OR4_680_Y), .C(OR4_452_Y), 
        .D(OR4_592_Y), .Y(R_DATA[0]));
    OR4 OR4_389 (.A(\R_DATA_TEMPR16[53] ), .B(\R_DATA_TEMPR17[53] ), 
        .C(\R_DATA_TEMPR18[53] ), .D(\R_DATA_TEMPR19[53] ), .Y(
        OR4_389_Y));
    OR4 OR4_392 (.A(OR4_474_Y), .B(OR4_231_Y), .C(OR4_478_Y), .D(
        OR4_215_Y), .Y(OR4_392_Y));
    OR4 OR4_19 (.A(OR4_147_Y), .B(OR4_576_Y), .C(OR4_0_Y), .D(
        OR4_363_Y), .Y(OR4_19_Y));
    OR4 OR4_41 (.A(\R_DATA_TEMPR16[49] ), .B(\R_DATA_TEMPR17[49] ), .C(
        \R_DATA_TEMPR18[49] ), .D(\R_DATA_TEMPR19[49] ), .Y(OR4_41_Y));
    OR4 OR4_333 (.A(\R_DATA_TEMPR16[63] ), .B(\R_DATA_TEMPR17[63] ), 
        .C(\R_DATA_TEMPR18[63] ), .D(\R_DATA_TEMPR19[63] ), .Y(
        OR4_333_Y));
    OR4 OR4_519 (.A(\R_DATA_TEMPR8[39] ), .B(\R_DATA_TEMPR9[39] ), .C(
        \R_DATA_TEMPR10[39] ), .D(\R_DATA_TEMPR11[39] ), .Y(OR4_519_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%17%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C1 (
        .A_DOUT({\R_DATA_TEMPR17[79] , \R_DATA_TEMPR17[78] , 
        \R_DATA_TEMPR17[77] , \R_DATA_TEMPR17[76] , 
        \R_DATA_TEMPR17[75] , \R_DATA_TEMPR17[74] , 
        \R_DATA_TEMPR17[73] , \R_DATA_TEMPR17[72] , 
        \R_DATA_TEMPR17[71] , \R_DATA_TEMPR17[70] , 
        \R_DATA_TEMPR17[69] , \R_DATA_TEMPR17[68] , 
        \R_DATA_TEMPR17[67] , \R_DATA_TEMPR17[66] , 
        \R_DATA_TEMPR17[65] , \R_DATA_TEMPR17[64] , 
        \R_DATA_TEMPR17[63] , \R_DATA_TEMPR17[62] , 
        \R_DATA_TEMPR17[61] , \R_DATA_TEMPR17[60] }), .B_DOUT({
        \R_DATA_TEMPR17[59] , \R_DATA_TEMPR17[58] , 
        \R_DATA_TEMPR17[57] , \R_DATA_TEMPR17[56] , 
        \R_DATA_TEMPR17[55] , \R_DATA_TEMPR17[54] , 
        \R_DATA_TEMPR17[53] , \R_DATA_TEMPR17[52] , 
        \R_DATA_TEMPR17[51] , \R_DATA_TEMPR17[50] , 
        \R_DATA_TEMPR17[49] , \R_DATA_TEMPR17[48] , 
        \R_DATA_TEMPR17[47] , \R_DATA_TEMPR17[46] , 
        \R_DATA_TEMPR17[45] , \R_DATA_TEMPR17[44] , 
        \R_DATA_TEMPR17[43] , \R_DATA_TEMPR17[42] , 
        \R_DATA_TEMPR17[41] , \R_DATA_TEMPR17[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[17][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_668 (.A(\R_DATA_TEMPR16[57] ), .B(\R_DATA_TEMPR17[57] ), 
        .C(\R_DATA_TEMPR18[57] ), .D(\R_DATA_TEMPR19[57] ), .Y(
        OR4_668_Y));
    OR4 OR4_510 (.A(\R_DATA_TEMPR24[46] ), .B(\R_DATA_TEMPR25[46] ), 
        .C(\R_DATA_TEMPR26[46] ), .D(\R_DATA_TEMPR27[46] ), .Y(
        OR4_510_Y));
    OR4 OR4_444 (.A(\R_DATA_TEMPR12[68] ), .B(\R_DATA_TEMPR13[68] ), 
        .C(\R_DATA_TEMPR14[68] ), .D(\R_DATA_TEMPR15[68] ), .Y(
        OR4_444_Y));
    OR4 OR4_432 (.A(\R_DATA_TEMPR0[78] ), .B(\R_DATA_TEMPR1[78] ), .C(
        \R_DATA_TEMPR2[78] ), .D(\R_DATA_TEMPR3[78] ), .Y(OR4_432_Y));
    OR4 OR4_528 (.A(\R_DATA_TEMPR8[13] ), .B(\R_DATA_TEMPR9[13] ), .C(
        \R_DATA_TEMPR10[13] ), .D(\R_DATA_TEMPR11[13] ), .Y(OR4_528_Y));
    OR2 OR2_76 (.A(\R_DATA_TEMPR20[13] ), .B(\R_DATA_TEMPR21[13] ), .Y(
        OR2_76_Y));
    OR4 OR4_52 (.A(\R_DATA_TEMPR8[56] ), .B(\R_DATA_TEMPR9[56] ), .C(
        \R_DATA_TEMPR10[56] ), .D(\R_DATA_TEMPR11[56] ), .Y(OR4_52_Y));
    OR4 OR4_662 (.A(OR4_432_Y), .B(OR4_289_Y), .C(OR4_169_Y), .D(
        OR4_220_Y), .Y(OR4_662_Y));
    OR4 OR4_439 (.A(OR4_15_Y), .B(OR4_267_Y), .C(OR4_566_Y), .D(
        OR4_134_Y), .Y(OR4_439_Y));
    OR4 OR4_346 (.A(\R_DATA_TEMPR8[54] ), .B(\R_DATA_TEMPR9[54] ), .C(
        \R_DATA_TEMPR10[54] ), .D(\R_DATA_TEMPR11[54] ), .Y(OR4_346_Y));
    OR4 OR4_136 (.A(OR4_56_Y), .B(OR2_62_Y), .C(\R_DATA_TEMPR22[4] ), 
        .D(\R_DATA_TEMPR23[4] ), .Y(OR4_136_Y));
    OR2 OR2_20 (.A(\R_DATA_TEMPR20[66] ), .B(\R_DATA_TEMPR21[66] ), .Y(
        OR2_20_Y));
    INV \INVBLKX1[0]  (.A(W_ADDR[10]), .Y(\BLKX1[0] ));
    OR2 OR2_16 (.A(\R_DATA_TEMPR20[48] ), .B(\R_DATA_TEMPR21[48] ), .Y(
        OR2_16_Y));
    CFG2 #( .INIT(4'h4) )  CFG2_6 (.A(R_ADDR[12]), .B(R_ADDR[11]), .Y(
        CFG2_6_Y));
    OR2 OR2_27 (.A(\R_DATA_TEMPR20[58] ), .B(\R_DATA_TEMPR21[58] ), .Y(
        OR2_27_Y));
    OR4 OR4_426 (.A(\R_DATA_TEMPR0[67] ), .B(\R_DATA_TEMPR1[67] ), .C(
        \R_DATA_TEMPR2[67] ), .D(\R_DATA_TEMPR3[67] ), .Y(OR4_426_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[0]  (.A(CFG2_3_Y), .B(
        R_ADDR[13]), .C(R_EN), .Y(\BLKY2[0] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%9%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0 (
        .A_DOUT({\R_DATA_TEMPR9[39] , \R_DATA_TEMPR9[38] , 
        \R_DATA_TEMPR9[37] , \R_DATA_TEMPR9[36] , \R_DATA_TEMPR9[35] , 
        \R_DATA_TEMPR9[34] , \R_DATA_TEMPR9[33] , \R_DATA_TEMPR9[32] , 
        \R_DATA_TEMPR9[31] , \R_DATA_TEMPR9[30] , \R_DATA_TEMPR9[29] , 
        \R_DATA_TEMPR9[28] , \R_DATA_TEMPR9[27] , \R_DATA_TEMPR9[26] , 
        \R_DATA_TEMPR9[25] , \R_DATA_TEMPR9[24] , \R_DATA_TEMPR9[23] , 
        \R_DATA_TEMPR9[22] , \R_DATA_TEMPR9[21] , \R_DATA_TEMPR9[20] })
        , .B_DOUT({\R_DATA_TEMPR9[19] , \R_DATA_TEMPR9[18] , 
        \R_DATA_TEMPR9[17] , \R_DATA_TEMPR9[16] , \R_DATA_TEMPR9[15] , 
        \R_DATA_TEMPR9[14] , \R_DATA_TEMPR9[13] , \R_DATA_TEMPR9[12] , 
        \R_DATA_TEMPR9[11] , \R_DATA_TEMPR9[10] , \R_DATA_TEMPR9[9] , 
        \R_DATA_TEMPR9[8] , \R_DATA_TEMPR9[7] , \R_DATA_TEMPR9[6] , 
        \R_DATA_TEMPR9[5] , \R_DATA_TEMPR9[4] , \R_DATA_TEMPR9[3] , 
        \R_DATA_TEMPR9[2] , \R_DATA_TEMPR9[1] , \R_DATA_TEMPR9[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[9][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_203 (.A(\R_DATA_TEMPR12[59] ), .B(\R_DATA_TEMPR13[59] ), 
        .C(\R_DATA_TEMPR14[59] ), .D(\R_DATA_TEMPR15[59] ), .Y(
        OR4_203_Y));
    OR4 OR4_290 (.A(\R_DATA_TEMPR24[59] ), .B(\R_DATA_TEMPR25[59] ), 
        .C(\R_DATA_TEMPR26[59] ), .D(\R_DATA_TEMPR27[59] ), .Y(
        OR4_290_Y));
    OR4 OR4_597 (.A(\R_DATA_TEMPR28[55] ), .B(\R_DATA_TEMPR29[55] ), 
        .C(\R_DATA_TEMPR30[55] ), .D(\R_DATA_TEMPR31[55] ), .Y(
        OR4_597_Y));
    OR4 OR4_338 (.A(OR4_111_Y), .B(OR4_694_Y), .C(OR4_574_Y), .D(
        OR4_609_Y), .Y(OR4_338_Y));
    OR4 OR4_273 (.A(\R_DATA_TEMPR4[47] ), .B(\R_DATA_TEMPR5[47] ), .C(
        \R_DATA_TEMPR6[47] ), .D(\R_DATA_TEMPR7[47] ), .Y(OR4_273_Y));
    OR4 \OR4_R_DATA[77]  (.A(OR4_117_Y), .B(OR4_473_Y), .C(OR4_657_Y), 
        .D(OR4_717_Y), .Y(R_DATA[77]));
    OR4 OR4_313 (.A(\R_DATA_TEMPR4[18] ), .B(\R_DATA_TEMPR5[18] ), .C(
        \R_DATA_TEMPR6[18] ), .D(\R_DATA_TEMPR7[18] ), .Y(OR4_313_Y));
    OR4 OR4_322 (.A(\R_DATA_TEMPR4[72] ), .B(\R_DATA_TEMPR5[72] ), .C(
        \R_DATA_TEMPR6[72] ), .D(\R_DATA_TEMPR7[72] ), .Y(OR4_322_Y));
    OR4 OR4_710 (.A(\R_DATA_TEMPR12[61] ), .B(\R_DATA_TEMPR13[61] ), 
        .C(\R_DATA_TEMPR14[61] ), .D(\R_DATA_TEMPR15[61] ), .Y(
        OR4_710_Y));
    OR4 OR4_699 (.A(\R_DATA_TEMPR4[74] ), .B(\R_DATA_TEMPR5[74] ), .C(
        \R_DATA_TEMPR6[74] ), .D(\R_DATA_TEMPR7[74] ), .Y(OR4_699_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%19%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0 (
        .A_DOUT({\R_DATA_TEMPR19[39] , \R_DATA_TEMPR19[38] , 
        \R_DATA_TEMPR19[37] , \R_DATA_TEMPR19[36] , 
        \R_DATA_TEMPR19[35] , \R_DATA_TEMPR19[34] , 
        \R_DATA_TEMPR19[33] , \R_DATA_TEMPR19[32] , 
        \R_DATA_TEMPR19[31] , \R_DATA_TEMPR19[30] , 
        \R_DATA_TEMPR19[29] , \R_DATA_TEMPR19[28] , 
        \R_DATA_TEMPR19[27] , \R_DATA_TEMPR19[26] , 
        \R_DATA_TEMPR19[25] , \R_DATA_TEMPR19[24] , 
        \R_DATA_TEMPR19[23] , \R_DATA_TEMPR19[22] , 
        \R_DATA_TEMPR19[21] , \R_DATA_TEMPR19[20] }), .B_DOUT({
        \R_DATA_TEMPR19[19] , \R_DATA_TEMPR19[18] , 
        \R_DATA_TEMPR19[17] , \R_DATA_TEMPR19[16] , 
        \R_DATA_TEMPR19[15] , \R_DATA_TEMPR19[14] , 
        \R_DATA_TEMPR19[13] , \R_DATA_TEMPR19[12] , 
        \R_DATA_TEMPR19[11] , \R_DATA_TEMPR19[10] , 
        \R_DATA_TEMPR19[9] , \R_DATA_TEMPR19[8] , \R_DATA_TEMPR19[7] , 
        \R_DATA_TEMPR19[6] , \R_DATA_TEMPR19[5] , \R_DATA_TEMPR19[4] , 
        \R_DATA_TEMPR19[3] , \R_DATA_TEMPR19[2] , \R_DATA_TEMPR19[1] , 
        \R_DATA_TEMPR19[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_12 (.A(\R_DATA_TEMPR0[58] ), .B(\R_DATA_TEMPR1[58] ), .C(
        \R_DATA_TEMPR2[58] ), .D(\R_DATA_TEMPR3[58] ), .Y(OR4_12_Y));
    OR4 OR4_583 (.A(\R_DATA_TEMPR4[75] ), .B(\R_DATA_TEMPR5[75] ), .C(
        \R_DATA_TEMPR6[75] ), .D(\R_DATA_TEMPR7[75] ), .Y(OR4_583_Y));
    OR4 OR4_412 (.A(OR4_654_Y), .B(OR4_507_Y), .C(OR4_498_Y), .D(
        OR4_227_Y), .Y(OR4_412_Y));
    OR4 OR4_296 (.A(\R_DATA_TEMPR12[49] ), .B(\R_DATA_TEMPR13[49] ), 
        .C(\R_DATA_TEMPR14[49] ), .D(\R_DATA_TEMPR15[49] ), .Y(
        OR4_296_Y));
    OR4 OR4_419 (.A(OR4_285_Y), .B(OR2_6_Y), .C(\R_DATA_TEMPR22[33] ), 
        .D(\R_DATA_TEMPR23[33] ), .Y(OR4_419_Y));
    OR4 OR4_251 (.A(\R_DATA_TEMPR16[55] ), .B(\R_DATA_TEMPR17[55] ), 
        .C(\R_DATA_TEMPR18[55] ), .D(\R_DATA_TEMPR19[55] ), .Y(
        OR4_251_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%11%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0 (
        .A_DOUT({\R_DATA_TEMPR11[39] , \R_DATA_TEMPR11[38] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR11[36] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR11[34] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR11[32] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR11[30] , 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR11[28] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR11[26] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR11[24] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR11[22] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR11[20] }), .B_DOUT({
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR11[18] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR11[16] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR11[14] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR11[12] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR11[10] , 
        \R_DATA_TEMPR11[9] , \R_DATA_TEMPR11[8] , \R_DATA_TEMPR11[7] , 
        \R_DATA_TEMPR11[6] , \R_DATA_TEMPR11[5] , \R_DATA_TEMPR11[4] , 
        \R_DATA_TEMPR11[3] , \R_DATA_TEMPR11[2] , \R_DATA_TEMPR11[1] , 
        \R_DATA_TEMPR11[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_79 (.A(\R_DATA_TEMPR8[50] ), .B(\R_DATA_TEMPR9[50] ), .C(
        \R_DATA_TEMPR10[50] ), .D(\R_DATA_TEMPR11[50] ), .Y(OR4_79_Y));
    OR4 OR4_139 (.A(\R_DATA_TEMPR28[23] ), .B(\R_DATA_TEMPR29[23] ), 
        .C(\R_DATA_TEMPR30[23] ), .D(\R_DATA_TEMPR31[23] ), .Y(
        OR4_139_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%14%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C1 (
        .A_DOUT({\R_DATA_TEMPR14[79] , \R_DATA_TEMPR14[78] , 
        \R_DATA_TEMPR14[77] , \R_DATA_TEMPR14[76] , 
        \R_DATA_TEMPR14[75] , \R_DATA_TEMPR14[74] , 
        \R_DATA_TEMPR14[73] , \R_DATA_TEMPR14[72] , 
        \R_DATA_TEMPR14[71] , \R_DATA_TEMPR14[70] , 
        \R_DATA_TEMPR14[69] , \R_DATA_TEMPR14[68] , 
        \R_DATA_TEMPR14[67] , \R_DATA_TEMPR14[66] , 
        \R_DATA_TEMPR14[65] , \R_DATA_TEMPR14[64] , 
        \R_DATA_TEMPR14[63] , \R_DATA_TEMPR14[62] , 
        \R_DATA_TEMPR14[61] , \R_DATA_TEMPR14[60] }), .B_DOUT({
        \R_DATA_TEMPR14[59] , \R_DATA_TEMPR14[58] , 
        \R_DATA_TEMPR14[57] , \R_DATA_TEMPR14[56] , 
        \R_DATA_TEMPR14[55] , \R_DATA_TEMPR14[54] , 
        \R_DATA_TEMPR14[53] , \R_DATA_TEMPR14[52] , 
        \R_DATA_TEMPR14[51] , \R_DATA_TEMPR14[50] , 
        \R_DATA_TEMPR14[49] , \R_DATA_TEMPR14[48] , 
        \R_DATA_TEMPR14[47] , \R_DATA_TEMPR14[46] , 
        \R_DATA_TEMPR14[45] , \R_DATA_TEMPR14[44] , 
        \R_DATA_TEMPR14[43] , \R_DATA_TEMPR14[42] , 
        \R_DATA_TEMPR14[41] , \R_DATA_TEMPR14[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[14][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[3] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_116 (.A(\R_DATA_TEMPR0[33] ), .B(\R_DATA_TEMPR1[33] ), .C(
        \R_DATA_TEMPR2[33] ), .D(\R_DATA_TEMPR3[33] ), .Y(OR4_116_Y));
    OR4 OR4_608 (.A(OR4_245_Y), .B(OR4_17_Y), .C(OR4_52_Y), .D(
        OR4_192_Y), .Y(OR4_608_Y));
    OR4 OR4_144 (.A(\R_DATA_TEMPR12[12] ), .B(\R_DATA_TEMPR13[12] ), 
        .C(\R_DATA_TEMPR14[12] ), .D(\R_DATA_TEMPR15[12] ), .Y(
        OR4_144_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%18%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0 (
        .A_DOUT({\R_DATA_TEMPR18[39] , \R_DATA_TEMPR18[38] , 
        \R_DATA_TEMPR18[37] , \R_DATA_TEMPR18[36] , 
        \R_DATA_TEMPR18[35] , \R_DATA_TEMPR18[34] , 
        \R_DATA_TEMPR18[33] , \R_DATA_TEMPR18[32] , 
        \R_DATA_TEMPR18[31] , \R_DATA_TEMPR18[30] , 
        \R_DATA_TEMPR18[29] , \R_DATA_TEMPR18[28] , 
        \R_DATA_TEMPR18[27] , \R_DATA_TEMPR18[26] , 
        \R_DATA_TEMPR18[25] , \R_DATA_TEMPR18[24] , 
        \R_DATA_TEMPR18[23] , \R_DATA_TEMPR18[22] , 
        \R_DATA_TEMPR18[21] , \R_DATA_TEMPR18[20] }), .B_DOUT({
        \R_DATA_TEMPR18[19] , \R_DATA_TEMPR18[18] , 
        \R_DATA_TEMPR18[17] , \R_DATA_TEMPR18[16] , 
        \R_DATA_TEMPR18[15] , \R_DATA_TEMPR18[14] , 
        \R_DATA_TEMPR18[13] , \R_DATA_TEMPR18[12] , 
        \R_DATA_TEMPR18[11] , \R_DATA_TEMPR18[10] , 
        \R_DATA_TEMPR18[9] , \R_DATA_TEMPR18[8] , \R_DATA_TEMPR18[7] , 
        \R_DATA_TEMPR18[6] , \R_DATA_TEMPR18[5] , \R_DATA_TEMPR18[4] , 
        \R_DATA_TEMPR18[3] , \R_DATA_TEMPR18[2] , \R_DATA_TEMPR18[1] , 
        \R_DATA_TEMPR18[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_694 (.A(\R_DATA_TEMPR4[48] ), .B(\R_DATA_TEMPR5[48] ), .C(
        \R_DATA_TEMPR6[48] ), .D(\R_DATA_TEMPR7[48] ), .Y(OR4_694_Y));
    OR2 OR2_70 (.A(\R_DATA_TEMPR20[43] ), .B(\R_DATA_TEMPR21[43] ), .Y(
        OR2_70_Y));
    OR4 OR4_678 (.A(\R_DATA_TEMPR12[37] ), .B(\R_DATA_TEMPR13[37] ), 
        .C(\R_DATA_TEMPR14[37] ), .D(\R_DATA_TEMPR15[37] ), .Y(
        OR4_678_Y));
    OR4 OR4_602 (.A(\R_DATA_TEMPR16[74] ), .B(\R_DATA_TEMPR17[74] ), 
        .C(\R_DATA_TEMPR18[74] ), .D(\R_DATA_TEMPR19[74] ), .Y(
        OR4_602_Y));
    OR4 \OR4_R_DATA[32]  (.A(OR4_690_Y), .B(OR4_672_Y), .C(OR4_567_Y), 
        .D(OR4_255_Y), .Y(R_DATA[32]));
    OR4 OR4_552 (.A(\R_DATA_TEMPR4[25] ), .B(\R_DATA_TEMPR5[25] ), .C(
        \R_DATA_TEMPR6[25] ), .D(\R_DATA_TEMPR7[25] ), .Y(OR4_552_Y));
    OR2 OR2_77 (.A(\R_DATA_TEMPR20[42] ), .B(\R_DATA_TEMPR21[42] ), .Y(
        OR2_77_Y));
    OR4 OR4_220 (.A(\R_DATA_TEMPR12[78] ), .B(\R_DATA_TEMPR13[78] ), 
        .C(\R_DATA_TEMPR14[78] ), .D(\R_DATA_TEMPR15[78] ), .Y(
        OR4_220_Y));
    OR4 OR4_672 (.A(OR4_360_Y), .B(OR2_14_Y), .C(\R_DATA_TEMPR22[32] ), 
        .D(\R_DATA_TEMPR23[32] ), .Y(OR4_672_Y));
    OR4 OR4_527 (.A(\R_DATA_TEMPR4[32] ), .B(\R_DATA_TEMPR5[32] ), .C(
        \R_DATA_TEMPR6[32] ), .D(\R_DATA_TEMPR7[32] ), .Y(OR4_527_Y));
    OR4 OR4_318 (.A(\R_DATA_TEMPR8[79] ), .B(\R_DATA_TEMPR9[79] ), .C(
        \R_DATA_TEMPR10[79] ), .D(\R_DATA_TEMPR11[79] ), .Y(OR4_318_Y));
    OR2 OR2_10 (.A(\R_DATA_TEMPR20[9] ), .B(\R_DATA_TEMPR21[9] ), .Y(
        OR2_10_Y));
    OR4 \OR4_R_DATA[55]  (.A(OR4_181_Y), .B(OR4_520_Y), .C(OR4_70_Y), 
        .D(OR4_597_Y), .Y(R_DATA[55]));
    OR4 \OR4_R_DATA[3]  (.A(OR4_178_Y), .B(OR4_373_Y), .C(OR4_314_Y), 
        .D(OR4_371_Y), .Y(R_DATA[3]));
    OR2 OR2_17 (.A(\R_DATA_TEMPR20[55] ), .B(\R_DATA_TEMPR21[55] ), .Y(
        OR2_17_Y));
    OR4 OR4_666 (.A(\R_DATA_TEMPR4[24] ), .B(\R_DATA_TEMPR5[24] ), .C(
        \R_DATA_TEMPR6[24] ), .D(\R_DATA_TEMPR7[24] ), .Y(OR4_666_Y));
    OR4 OR4_629 (.A(\R_DATA_TEMPR0[26] ), .B(\R_DATA_TEMPR1[26] ), .C(
        \R_DATA_TEMPR2[26] ), .D(\R_DATA_TEMPR3[26] ), .Y(OR4_629_Y));
    OR4 OR4_554 (.A(\R_DATA_TEMPR4[27] ), .B(\R_DATA_TEMPR5[27] ), .C(
        \R_DATA_TEMPR6[27] ), .D(\R_DATA_TEMPR7[27] ), .Y(OR4_554_Y));
    OR4 OR4_546 (.A(\R_DATA_TEMPR28[65] ), .B(\R_DATA_TEMPR29[65] ), 
        .C(\R_DATA_TEMPR30[65] ), .D(\R_DATA_TEMPR31[65] ), .Y(
        OR4_546_Y));
    OR4 OR4_226 (.A(\R_DATA_TEMPR4[64] ), .B(\R_DATA_TEMPR5[64] ), .C(
        \R_DATA_TEMPR6[64] ), .D(\R_DATA_TEMPR7[64] ), .Y(OR4_226_Y));
    OR4 OR4_119 (.A(\R_DATA_TEMPR24[37] ), .B(\R_DATA_TEMPR25[37] ), 
        .C(\R_DATA_TEMPR26[37] ), .D(\R_DATA_TEMPR27[37] ), .Y(
        OR4_119_Y));
    OR4 OR4_72 (.A(\R_DATA_TEMPR0[50] ), .B(\R_DATA_TEMPR1[50] ), .C(
        \R_DATA_TEMPR2[50] ), .D(\R_DATA_TEMPR3[50] ), .Y(OR4_72_Y));
    OR4 OR4_637 (.A(\R_DATA_TEMPR16[25] ), .B(\R_DATA_TEMPR17[25] ), 
        .C(\R_DATA_TEMPR18[25] ), .D(\R_DATA_TEMPR19[25] ), .Y(
        OR4_637_Y));
    OR4 OR4_624 (.A(\R_DATA_TEMPR24[27] ), .B(\R_DATA_TEMPR25[27] ), 
        .C(\R_DATA_TEMPR26[27] ), .D(\R_DATA_TEMPR27[27] ), .Y(
        OR4_624_Y));
    OR4 OR4_351 (.A(\R_DATA_TEMPR4[70] ), .B(\R_DATA_TEMPR5[70] ), .C(
        \R_DATA_TEMPR6[70] ), .D(\R_DATA_TEMPR7[70] ), .Y(OR4_351_Y));
    OR2 OR2_28 (.A(\R_DATA_TEMPR20[14] ), .B(\R_DATA_TEMPR21[14] ), .Y(
        OR2_28_Y));
    OR4 \OR4_R_DATA[33]  (.A(OR4_611_Y), .B(OR4_419_Y), .C(OR4_391_Y), 
        .D(OR4_366_Y), .Y(R_DATA[33]));
    OR4 OR4_450 (.A(\R_DATA_TEMPR12[27] ), .B(\R_DATA_TEMPR13[27] ), 
        .C(\R_DATA_TEMPR14[27] ), .D(\R_DATA_TEMPR15[27] ), .Y(
        OR4_450_Y));
    OR4 \OR4_R_DATA[25]  (.A(OR4_571_Y), .B(OR4_205_Y), .C(OR4_472_Y), 
        .D(OR4_274_Y), .Y(R_DATA[25]));
    OR4 OR4_283 (.A(\R_DATA_TEMPR24[64] ), .B(\R_DATA_TEMPR25[64] ), 
        .C(\R_DATA_TEMPR26[64] ), .D(\R_DATA_TEMPR27[64] ), .Y(
        OR4_283_Y));
    OR4 OR4_96 (.A(\R_DATA_TEMPR4[7] ), .B(\R_DATA_TEMPR5[7] ), .C(
        \R_DATA_TEMPR6[7] ), .D(\R_DATA_TEMPR7[7] ), .Y(OR4_96_Y));
    OR4 OR4_548 (.A(\R_DATA_TEMPR28[46] ), .B(\R_DATA_TEMPR29[46] ), 
        .C(\R_DATA_TEMPR30[46] ), .D(\R_DATA_TEMPR31[46] ), .Y(
        OR4_548_Y));
    OR4 OR4_54 (.A(\R_DATA_TEMPR28[70] ), .B(\R_DATA_TEMPR29[70] ), .C(
        \R_DATA_TEMPR30[70] ), .D(\R_DATA_TEMPR31[70] ), .Y(OR4_54_Y));
    OR4 OR4_3 (.A(OR4_102_Y), .B(OR2_72_Y), .C(\R_DATA_TEMPR22[70] ), 
        .D(\R_DATA_TEMPR23[70] ), .Y(OR4_3_Y));
    OR4 OR4_364 (.A(\R_DATA_TEMPR12[60] ), .B(\R_DATA_TEMPR13[60] ), 
        .C(\R_DATA_TEMPR14[60] ), .D(\R_DATA_TEMPR15[60] ), .Y(
        OR4_364_Y));
    OR4 OR4_606 (.A(\R_DATA_TEMPR16[69] ), .B(\R_DATA_TEMPR17[69] ), 
        .C(\R_DATA_TEMPR18[69] ), .D(\R_DATA_TEMPR19[69] ), .Y(
        OR4_606_Y));
    OR4 OR4_715 (.A(OR4_616_Y), .B(OR2_78_Y), .C(\R_DATA_TEMPR22[67] ), 
        .D(\R_DATA_TEMPR23[67] ), .Y(OR4_715_Y));
    OR4 OR4_617 (.A(\R_DATA_TEMPR12[79] ), .B(\R_DATA_TEMPR13[79] ), 
        .C(\R_DATA_TEMPR14[79] ), .D(\R_DATA_TEMPR15[79] ), .Y(
        OR4_617_Y));
    OR4 OR4_446 (.A(\R_DATA_TEMPR8[26] ), .B(\R_DATA_TEMPR9[26] ), .C(
        \R_DATA_TEMPR10[26] ), .D(\R_DATA_TEMPR11[26] ), .Y(OR4_446_Y));
    OR4 OR4_161 (.A(\R_DATA_TEMPR0[75] ), .B(\R_DATA_TEMPR1[75] ), .C(
        \R_DATA_TEMPR2[75] ), .D(\R_DATA_TEMPR3[75] ), .Y(OR4_161_Y));
    OR4 OR4_716 (.A(OR4_408_Y), .B(OR2_41_Y), .C(\R_DATA_TEMPR22[62] ), 
        .D(\R_DATA_TEMPR23[62] ), .Y(OR4_716_Y));
    OR4 OR4_676 (.A(\R_DATA_TEMPR8[36] ), .B(\R_DATA_TEMPR9[36] ), .C(
        \R_DATA_TEMPR10[36] ), .D(\R_DATA_TEMPR11[36] ), .Y(OR4_676_Y));
    OR4 OR4_237 (.A(\R_DATA_TEMPR12[25] ), .B(\R_DATA_TEMPR13[25] ), 
        .C(\R_DATA_TEMPR14[25] ), .D(\R_DATA_TEMPR15[25] ), .Y(
        OR4_237_Y));
    OR4 OR4_688 (.A(OR4_105_Y), .B(OR2_13_Y), .C(\R_DATA_TEMPR22[5] ), 
        .D(\R_DATA_TEMPR23[5] ), .Y(OR4_688_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%23%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0 (
        .A_DOUT({\R_DATA_TEMPR23[39] , \R_DATA_TEMPR23[38] , 
        \R_DATA_TEMPR23[37] , \R_DATA_TEMPR23[36] , 
        \R_DATA_TEMPR23[35] , \R_DATA_TEMPR23[34] , 
        \R_DATA_TEMPR23[33] , \R_DATA_TEMPR23[32] , 
        \R_DATA_TEMPR23[31] , \R_DATA_TEMPR23[30] , 
        \R_DATA_TEMPR23[29] , \R_DATA_TEMPR23[28] , 
        \R_DATA_TEMPR23[27] , \R_DATA_TEMPR23[26] , 
        \R_DATA_TEMPR23[25] , \R_DATA_TEMPR23[24] , 
        \R_DATA_TEMPR23[23] , \R_DATA_TEMPR23[22] , 
        \R_DATA_TEMPR23[21] , \R_DATA_TEMPR23[20] }), .B_DOUT({
        \R_DATA_TEMPR23[19] , \R_DATA_TEMPR23[18] , 
        \R_DATA_TEMPR23[17] , \R_DATA_TEMPR23[16] , 
        \R_DATA_TEMPR23[15] , \R_DATA_TEMPR23[14] , 
        \R_DATA_TEMPR23[13] , \R_DATA_TEMPR23[12] , 
        \R_DATA_TEMPR23[11] , \R_DATA_TEMPR23[10] , 
        \R_DATA_TEMPR23[9] , \R_DATA_TEMPR23[8] , \R_DATA_TEMPR23[7] , 
        \R_DATA_TEMPR23[6] , \R_DATA_TEMPR23[5] , \R_DATA_TEMPR23[4] , 
        \R_DATA_TEMPR23[3] , \R_DATA_TEMPR23[2] , \R_DATA_TEMPR23[1] , 
        \R_DATA_TEMPR23[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_137 (.A(\R_DATA_TEMPR8[77] ), .B(\R_DATA_TEMPR9[77] ), .C(
        \R_DATA_TEMPR10[77] ), .D(\R_DATA_TEMPR11[77] ), .Y(OR4_137_Y));
    OR2 OR2_78 (.A(\R_DATA_TEMPR20[67] ), .B(\R_DATA_TEMPR21[67] ), .Y(
        OR2_78_Y));
    OR4 OR4_682 (.A(\R_DATA_TEMPR24[17] ), .B(\R_DATA_TEMPR25[17] ), 
        .C(\R_DATA_TEMPR26[17] ), .D(\R_DATA_TEMPR27[17] ), .Y(
        OR4_682_Y));
    OR4 OR4_342 (.A(\R_DATA_TEMPR4[71] ), .B(\R_DATA_TEMPR5[71] ), .C(
        \R_DATA_TEMPR6[71] ), .D(\R_DATA_TEMPR7[71] ), .Y(OR4_342_Y));
    OR4 OR4_461 (.A(\R_DATA_TEMPR16[52] ), .B(\R_DATA_TEMPR17[52] ), 
        .C(\R_DATA_TEMPR18[52] ), .D(\R_DATA_TEMPR19[52] ), .Y(
        OR4_461_Y));
    OR4 OR4_359 (.A(\R_DATA_TEMPR24[10] ), .B(\R_DATA_TEMPR25[10] ), 
        .C(\R_DATA_TEMPR26[10] ), .D(\R_DATA_TEMPR27[10] ), .Y(
        OR4_359_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%6%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C1 (
        .A_DOUT({\R_DATA_TEMPR6[79] , \R_DATA_TEMPR6[78] , 
        \R_DATA_TEMPR6[77] , \R_DATA_TEMPR6[76] , \R_DATA_TEMPR6[75] , 
        \R_DATA_TEMPR6[74] , \R_DATA_TEMPR6[73] , \R_DATA_TEMPR6[72] , 
        \R_DATA_TEMPR6[71] , \R_DATA_TEMPR6[70] , \R_DATA_TEMPR6[69] , 
        \R_DATA_TEMPR6[68] , \R_DATA_TEMPR6[67] , \R_DATA_TEMPR6[66] , 
        \R_DATA_TEMPR6[65] , \R_DATA_TEMPR6[64] , \R_DATA_TEMPR6[63] , 
        \R_DATA_TEMPR6[62] , \R_DATA_TEMPR6[61] , \R_DATA_TEMPR6[60] })
        , .B_DOUT({\R_DATA_TEMPR6[59] , \R_DATA_TEMPR6[58] , 
        \R_DATA_TEMPR6[57] , \R_DATA_TEMPR6[56] , \R_DATA_TEMPR6[55] , 
        \R_DATA_TEMPR6[54] , \R_DATA_TEMPR6[53] , \R_DATA_TEMPR6[52] , 
        \R_DATA_TEMPR6[51] , \R_DATA_TEMPR6[50] , \R_DATA_TEMPR6[49] , 
        \R_DATA_TEMPR6[48] , \R_DATA_TEMPR6[47] , \R_DATA_TEMPR6[46] , 
        \R_DATA_TEMPR6[45] , \R_DATA_TEMPR6[44] , \R_DATA_TEMPR6[43] , 
        \R_DATA_TEMPR6[42] , \R_DATA_TEMPR6[41] , \R_DATA_TEMPR6[40] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[6][1] ), .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], 
        R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], 
        R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({\BLKY2[1] , 
        R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA[79], 
        W_DATA[78], W_DATA[77], W_DATA[76], W_DATA[75], W_DATA[74], 
        W_DATA[73], W_DATA[72], W_DATA[71], W_DATA[70], W_DATA[69], 
        W_DATA[68], W_DATA[67], W_DATA[66], W_DATA[65], W_DATA[64], 
        W_DATA[63], W_DATA[62], W_DATA[61], W_DATA[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, GND}), 
        .B_BLK_EN({\BLKX2[1] , W_ADDR[10], \BLKX0[0] }), .B_CLK(CLK), 
        .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_14 (.A(\R_DATA_TEMPR0[34] ), .B(\R_DATA_TEMPR1[34] ), .C(
        \R_DATA_TEMPR2[34] ), .D(\R_DATA_TEMPR3[34] ), .Y(OR4_14_Y));
    OR4 OR4_468 (.A(OR4_198_Y), .B(OR2_53_Y), .C(\R_DATA_TEMPR22[65] ), 
        .D(\R_DATA_TEMPR23[65] ), .Y(OR4_468_Y));
    OR2 OR2_18 (.A(\R_DATA_TEMPR20[15] ), .B(\R_DATA_TEMPR21[15] ), .Y(
        OR2_18_Y));
    OR4 OR4_291 (.A(\R_DATA_TEMPR8[45] ), .B(\R_DATA_TEMPR9[45] ), .C(
        \R_DATA_TEMPR10[45] ), .D(\R_DATA_TEMPR11[45] ), .Y(OR4_291_Y));
    OR4 OR4_234 (.A(OR4_667_Y), .B(OR2_73_Y), .C(\R_DATA_TEMPR22[75] ), 
        .D(\R_DATA_TEMPR23[75] ), .Y(OR4_234_Y));
    OR4 OR4_90 (.A(OR4_239_Y), .B(OR4_639_Y), .C(OR4_399_Y), .D(
        OR4_157_Y), .Y(OR4_90_Y));
    OR4 OR4_46 (.A(\R_DATA_TEMPR16[47] ), .B(\R_DATA_TEMPR17[47] ), .C(
        \R_DATA_TEMPR18[47] ), .D(\R_DATA_TEMPR19[47] ), .Y(OR4_46_Y));
    OR4 OR4_569 (.A(\R_DATA_TEMPR16[24] ), .B(\R_DATA_TEMPR17[24] ), 
        .C(\R_DATA_TEMPR18[24] ), .D(\R_DATA_TEMPR19[24] ), .Y(
        OR4_569_Y));
    OR4 OR4_97 (.A(\R_DATA_TEMPR24[76] ), .B(\R_DATA_TEMPR25[76] ), .C(
        \R_DATA_TEMPR26[76] ), .D(\R_DATA_TEMPR27[76] ), .Y(OR4_97_Y));
    OR4 \OR4_R_DATA[6]  (.A(OR4_168_Y), .B(OR4_515_Y), .C(OR4_27_Y), 
        .D(OR4_118_Y), .Y(R_DATA[6]));
    OR4 OR4_592 (.A(\R_DATA_TEMPR28[0] ), .B(\R_DATA_TEMPR29[0] ), .C(
        \R_DATA_TEMPR30[0] ), .D(\R_DATA_TEMPR31[0] ), .Y(OR4_592_Y));
    OR4 OR4_63 (.A(\R_DATA_TEMPR8[1] ), .B(\R_DATA_TEMPR9[1] ), .C(
        \R_DATA_TEMPR10[1] ), .D(\R_DATA_TEMPR11[1] ), .Y(OR4_63_Y));
    OR4 OR4_560 (.A(\R_DATA_TEMPR28[9] ), .B(\R_DATA_TEMPR29[9] ), .C(
        \R_DATA_TEMPR30[9] ), .D(\R_DATA_TEMPR31[9] ), .Y(OR4_560_Y));
    OR4 OR4_217 (.A(\R_DATA_TEMPR24[28] ), .B(\R_DATA_TEMPR25[28] ), 
        .C(\R_DATA_TEMPR26[28] ), .D(\R_DATA_TEMPR27[28] ), .Y(
        OR4_217_Y));
    OR4 OR4_240 (.A(OR4_524_Y), .B(OR4_40_Y), .C(OR4_347_Y), .D(
        OR4_649_Y), .Y(OR4_240_Y));
    OR4 OR4_304 (.A(\R_DATA_TEMPR4[59] ), .B(\R_DATA_TEMPR5[59] ), .C(
        \R_DATA_TEMPR6[59] ), .D(\R_DATA_TEMPR7[59] ), .Y(OR4_304_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%20%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C1 (
        .A_DOUT({\R_DATA_TEMPR20[79] , \R_DATA_TEMPR20[78] , 
        \R_DATA_TEMPR20[77] , \R_DATA_TEMPR20[76] , 
        \R_DATA_TEMPR20[75] , \R_DATA_TEMPR20[74] , 
        \R_DATA_TEMPR20[73] , \R_DATA_TEMPR20[72] , 
        \R_DATA_TEMPR20[71] , \R_DATA_TEMPR20[70] , 
        \R_DATA_TEMPR20[69] , \R_DATA_TEMPR20[68] , 
        \R_DATA_TEMPR20[67] , \R_DATA_TEMPR20[66] , 
        \R_DATA_TEMPR20[65] , \R_DATA_TEMPR20[64] , 
        \R_DATA_TEMPR20[63] , \R_DATA_TEMPR20[62] , 
        \R_DATA_TEMPR20[61] , \R_DATA_TEMPR20[60] }), .B_DOUT({
        \R_DATA_TEMPR20[59] , \R_DATA_TEMPR20[58] , 
        \R_DATA_TEMPR20[57] , \R_DATA_TEMPR20[56] , 
        \R_DATA_TEMPR20[55] , \R_DATA_TEMPR20[54] , 
        \R_DATA_TEMPR20[53] , \R_DATA_TEMPR20[52] , 
        \R_DATA_TEMPR20[51] , \R_DATA_TEMPR20[50] , 
        \R_DATA_TEMPR20[49] , \R_DATA_TEMPR20[48] , 
        \R_DATA_TEMPR20[47] , \R_DATA_TEMPR20[46] , 
        \R_DATA_TEMPR20[45] , \R_DATA_TEMPR20[44] , 
        \R_DATA_TEMPR20[43] , \R_DATA_TEMPR20[42] , 
        \R_DATA_TEMPR20[41] , \R_DATA_TEMPR20[40] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[20][1] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[79], W_DATA[78], W_DATA[77], W_DATA[76], 
        W_DATA[75], W_DATA[74], W_DATA[73], W_DATA[72], W_DATA[71], 
        W_DATA[70], W_DATA[69], W_DATA[68], W_DATA[67], W_DATA[66], 
        W_DATA[65], W_DATA[64], W_DATA[63], W_DATA[62], W_DATA[61], 
        W_DATA[60]}), .A_REN(VCC), .A_WEN({WBYTE_EN[7], WBYTE_EN[6]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[59], W_DATA[58], W_DATA[57], W_DATA[56], 
        W_DATA[55], W_DATA[54], W_DATA[53], W_DATA[52], W_DATA[51], 
        W_DATA[50], W_DATA[49], W_DATA[48], W_DATA[47], W_DATA[46], 
        W_DATA[45], W_DATA[44], W_DATA[43], W_DATA[42], W_DATA[41], 
        W_DATA[40]}), .B_REN(VCC), .B_WEN({WBYTE_EN[5], WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_117 (.A(OR4_195_Y), .B(OR4_584_Y), .C(OR4_137_Y), .D(
        OR4_489_Y), .Y(OR4_117_Y));
    OR4 OR4_547 (.A(\R_DATA_TEMPR28[34] ), .B(\R_DATA_TEMPR29[34] ), 
        .C(\R_DATA_TEMPR30[34] ), .D(\R_DATA_TEMPR31[34] ), .Y(
        OR4_547_Y));
    OR4 OR4_335 (.A(OR4_232_Y), .B(OR4_376_Y), .C(OR4_451_Y), .D(
        OR4_270_Y), .Y(OR4_335_Y));
    OR4 OR4_374 (.A(OR4_569_Y), .B(OR2_51_Y), .C(\R_DATA_TEMPR22[24] ), 
        .D(\R_DATA_TEMPR23[24] ), .Y(OR4_374_Y));
    OR4 \OR4_R_DATA[1]  (.A(OR4_589_Y), .B(OR4_677_Y), .C(OR4_480_Y), 
        .D(OR4_384_Y), .Y(R_DATA[1]));
    OR4 OR4_101 (.A(\R_DATA_TEMPR28[26] ), .B(\R_DATA_TEMPR29[26] ), 
        .C(\R_DATA_TEMPR30[26] ), .D(\R_DATA_TEMPR31[26] ), .Y(
        OR4_101_Y));
    OR4 OR4_649 (.A(\R_DATA_TEMPR12[19] ), .B(\R_DATA_TEMPR13[19] ), 
        .C(\R_DATA_TEMPR14[19] ), .D(\R_DATA_TEMPR15[19] ), .Y(
        OR4_649_Y));
    OR4 OR4_594 (.A(OR4_222_Y), .B(OR2_29_Y), .C(\R_DATA_TEMPR22[18] ), 
        .D(\R_DATA_TEMPR23[18] ), .Y(OR4_594_Y));
    OR4 OR4_171 (.A(OR4_458_Y), .B(OR4_704_Y), .C(OR4_288_Y), .D(
        OR4_585_Y), .Y(OR4_171_Y));
    OR4 OR4_713 (.A(OR4_334_Y), .B(OR4_114_Y), .C(OR4_160_Y), .D(
        OR4_287_Y), .Y(OR4_713_Y));
    OR4 OR4_553 (.A(\R_DATA_TEMPR16[46] ), .B(\R_DATA_TEMPR17[46] ), 
        .C(\R_DATA_TEMPR18[46] ), .D(\R_DATA_TEMPR19[46] ), .Y(
        OR4_553_Y));
    OR4 OR4_214 (.A(OR4_306_Y), .B(OR2_25_Y), .C(\R_DATA_TEMPR22[30] ), 
        .D(\R_DATA_TEMPR23[30] ), .Y(OR4_214_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%10%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0 (
        .A_DOUT({\R_DATA_TEMPR10[39] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR10[37] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR10[35] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR10[33] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR10[31] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR10[29] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR10[27] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR10[25] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR10[23] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR10[21] , \R_DATA_TEMPR10[20] }), .B_DOUT({
        \R_DATA_TEMPR10[19] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR10[17] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR10[15] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR10[13] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR10[11] , \R_DATA_TEMPR10[10] , 
        \R_DATA_TEMPR10[9] , \R_DATA_TEMPR10[8] , \R_DATA_TEMPR10[7] , 
        \R_DATA_TEMPR10[6] , \R_DATA_TEMPR10[5] , \R_DATA_TEMPR10[4] , 
        \R_DATA_TEMPR10[3] , \R_DATA_TEMPR10[2] , \R_DATA_TEMPR10[1] , 
        \R_DATA_TEMPR10[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_246 (.A(\R_DATA_TEMPR24[4] ), .B(\R_DATA_TEMPR25[4] ), .C(
        \R_DATA_TEMPR26[4] ), .D(\R_DATA_TEMPR27[4] ), .Y(OR4_246_Y));
    OR4 OR4_221 (.A(\R_DATA_TEMPR4[39] ), .B(\R_DATA_TEMPR5[39] ), .C(
        \R_DATA_TEMPR6[39] ), .D(\R_DATA_TEMPR7[39] ), .Y(OR4_221_Y));
    OR4 OR4_401 (.A(\R_DATA_TEMPR24[56] ), .B(\R_DATA_TEMPR25[56] ), 
        .C(\R_DATA_TEMPR26[56] ), .D(\R_DATA_TEMPR27[56] ), .Y(
        OR4_401_Y));
    OR4 \OR4_R_DATA[58]  (.A(OR4_249_Y), .B(OR4_133_Y), .C(OR4_532_Y), 
        .D(OR4_634_Y), .Y(R_DATA[58]));
    OR4 OR4_74 (.A(\R_DATA_TEMPR16[20] ), .B(\R_DATA_TEMPR17[20] ), .C(
        \R_DATA_TEMPR18[20] ), .D(\R_DATA_TEMPR19[20] ), .Y(OR4_74_Y));
    OR4 OR4_408 (.A(\R_DATA_TEMPR16[62] ), .B(\R_DATA_TEMPR17[62] ), 
        .C(\R_DATA_TEMPR18[62] ), .D(\R_DATA_TEMPR19[62] ), .Y(
        OR4_408_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[6]  (.A(CFG2_7_Y), .B(
        W_ADDR[13]), .C(W_EN), .Y(\BLKX2[6] ));
    OR4 OR4_471 (.A(\R_DATA_TEMPR4[16] ), .B(\R_DATA_TEMPR5[16] ), .C(
        \R_DATA_TEMPR6[16] ), .D(\R_DATA_TEMPR7[16] ), .Y(OR4_471_Y));
    OR4 OR4_363 (.A(\R_DATA_TEMPR12[62] ), .B(\R_DATA_TEMPR13[62] ), 
        .C(\R_DATA_TEMPR14[62] ), .D(\R_DATA_TEMPR15[62] ), .Y(
        OR4_363_Y));
    OR4 OR4_478 (.A(\R_DATA_TEMPR8[2] ), .B(\R_DATA_TEMPR9[2] ), .C(
        \R_DATA_TEMPR10[2] ), .D(\R_DATA_TEMPR11[2] ), .Y(OR4_478_Y));
    OR4 OR4_391 (.A(\R_DATA_TEMPR24[33] ), .B(\R_DATA_TEMPR25[33] ), 
        .C(\R_DATA_TEMPR26[33] ), .D(\R_DATA_TEMPR27[33] ), .Y(
        OR4_391_Y));
    OR4 OR4_644 (.A(\R_DATA_TEMPR4[36] ), .B(\R_DATA_TEMPR5[36] ), .C(
        \R_DATA_TEMPR6[36] ), .D(\R_DATA_TEMPR7[36] ), .Y(OR4_644_Y));
    OR4 OR4_61 (.A(\R_DATA_TEMPR0[59] ), .B(\R_DATA_TEMPR1[59] ), .C(
        \R_DATA_TEMPR2[59] ), .D(\R_DATA_TEMPR3[59] ), .Y(OR4_61_Y));
    OR4 OR4_462 (.A(OR4_596_Y), .B(OR4_297_Y), .C(OR4_445_Y), .D(
        OR4_80_Y), .Y(OR4_462_Y));
    OR4 OR4_635 (.A(OR4_110_Y), .B(OR2_56_Y), .C(\R_DATA_TEMPR22[21] ), 
        .D(\R_DATA_TEMPR23[21] ), .Y(OR4_635_Y));
    OR4 OR4_522 (.A(\R_DATA_TEMPR12[42] ), .B(\R_DATA_TEMPR13[42] ), 
        .C(\R_DATA_TEMPR14[42] ), .D(\R_DATA_TEMPR15[42] ), .Y(
        OR4_522_Y));
    OR4 OR4_686 (.A(OR4_572_Y), .B(OR4_718_Y), .C(OR4_71_Y), .D(
        OR4_610_Y), .Y(OR4_686_Y));
    OR4 OR4_469 (.A(OR4_333_Y), .B(OR2_34_Y), .C(\R_DATA_TEMPR22[63] ), 
        .D(\R_DATA_TEMPR23[63] ), .Y(OR4_469_Y));
    OR2 OR2_5 (.A(\R_DATA_TEMPR20[40] ), .B(\R_DATA_TEMPR21[40] ), .Y(
        OR2_5_Y));
    OR4 OR4_315 (.A(\R_DATA_TEMPR28[24] ), .B(\R_DATA_TEMPR29[24] ), 
        .C(\R_DATA_TEMPR30[24] ), .D(\R_DATA_TEMPR31[24] ), .Y(
        OR4_315_Y));
    OR4 OR4_490 (.A(\R_DATA_TEMPR16[2] ), .B(\R_DATA_TEMPR17[2] ), .C(
        \R_DATA_TEMPR18[2] ), .D(\R_DATA_TEMPR19[2] ), .Y(OR4_490_Y));
    OR4 OR4_40 (.A(\R_DATA_TEMPR4[19] ), .B(\R_DATA_TEMPR5[19] ), .C(
        \R_DATA_TEMPR6[19] ), .D(\R_DATA_TEMPR7[19] ), .Y(OR4_40_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%5%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0 (
        .A_DOUT({\R_DATA_TEMPR5[39] , \R_DATA_TEMPR5[38] , 
        \R_DATA_TEMPR5[37] , \R_DATA_TEMPR5[36] , \R_DATA_TEMPR5[35] , 
        \R_DATA_TEMPR5[34] , \R_DATA_TEMPR5[33] , \R_DATA_TEMPR5[32] , 
        \R_DATA_TEMPR5[31] , \R_DATA_TEMPR5[30] , \R_DATA_TEMPR5[29] , 
        \R_DATA_TEMPR5[28] , \R_DATA_TEMPR5[27] , \R_DATA_TEMPR5[26] , 
        \R_DATA_TEMPR5[25] , \R_DATA_TEMPR5[24] , \R_DATA_TEMPR5[23] , 
        \R_DATA_TEMPR5[22] , \R_DATA_TEMPR5[21] , \R_DATA_TEMPR5[20] })
        , .B_DOUT({\R_DATA_TEMPR5[19] , \R_DATA_TEMPR5[18] , 
        \R_DATA_TEMPR5[17] , \R_DATA_TEMPR5[16] , \R_DATA_TEMPR5[15] , 
        \R_DATA_TEMPR5[14] , \R_DATA_TEMPR5[13] , \R_DATA_TEMPR5[12] , 
        \R_DATA_TEMPR5[11] , \R_DATA_TEMPR5[10] , \R_DATA_TEMPR5[9] , 
        \R_DATA_TEMPR5[8] , \R_DATA_TEMPR5[7] , \R_DATA_TEMPR5[6] , 
        \R_DATA_TEMPR5[5] , \R_DATA_TEMPR5[4] , \R_DATA_TEMPR5[3] , 
        \R_DATA_TEMPR5[2] , \R_DATA_TEMPR5[1] , \R_DATA_TEMPR5[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[5][0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_509 (.A(\R_DATA_TEMPR8[16] ), .B(\R_DATA_TEMPR9[16] ), .C(
        \R_DATA_TEMPR10[16] ), .D(\R_DATA_TEMPR11[16] ), .Y(OR4_509_Y));
    OR4 OR4_166 (.A(\R_DATA_TEMPR4[34] ), .B(\R_DATA_TEMPR5[34] ), .C(
        \R_DATA_TEMPR6[34] ), .D(\R_DATA_TEMPR7[34] ), .Y(OR4_166_Y));
    OR4 OR4_500 (.A(\R_DATA_TEMPR12[58] ), .B(\R_DATA_TEMPR13[58] ), 
        .C(\R_DATA_TEMPR14[58] ), .D(\R_DATA_TEMPR15[58] ), .Y(
        OR4_500_Y));
    OR4 OR4_47 (.A(\R_DATA_TEMPR12[34] ), .B(\R_DATA_TEMPR13[34] ), .C(
        \R_DATA_TEMPR14[34] ), .D(\R_DATA_TEMPR15[34] ), .Y(OR4_47_Y));
    OR4 OR4_579 (.A(\R_DATA_TEMPR12[26] ), .B(\R_DATA_TEMPR13[26] ), 
        .C(\R_DATA_TEMPR14[26] ), .D(\R_DATA_TEMPR15[26] ), .Y(
        OR4_579_Y));
    OR4 OR4_570 (.A(\R_DATA_TEMPR16[42] ), .B(\R_DATA_TEMPR17[42] ), 
        .C(\R_DATA_TEMPR18[42] ), .D(\R_DATA_TEMPR19[42] ), .Y(
        OR4_570_Y));
    OR4 OR4_524 (.A(\R_DATA_TEMPR0[19] ), .B(\R_DATA_TEMPR1[19] ), .C(
        \R_DATA_TEMPR2[19] ), .D(\R_DATA_TEMPR3[19] ), .Y(OR4_524_Y));
    OR4 \OR4_R_DATA[28]  (.A(OR4_633_Y), .B(OR4_536_Y), .C(OR4_217_Y), 
        .D(OR4_303_Y), .Y(R_DATA[28]));
    OR4 OR4_368 (.A(\R_DATA_TEMPR4[11] ), .B(\R_DATA_TEMPR5[11] ), .C(
        \R_DATA_TEMPR6[11] ), .D(\R_DATA_TEMPR7[11] ), .Y(OR4_368_Y));
    OR4 OR4_712 (.A(OR4_238_Y), .B(OR4_75_Y), .C(OR4_64_Y), .D(
        OR4_514_Y), .Y(OR4_712_Y));
    OR4 OR4_630 (.A(OR4_511_Y), .B(OR4_666_Y), .C(OR4_20_Y), .D(
        OR4_550_Y), .Y(OR4_630_Y));
    OR4 OR4_98 (.A(\R_DATA_TEMPR8[27] ), .B(\R_DATA_TEMPR9[27] ), .C(
        \R_DATA_TEMPR10[27] ), .D(\R_DATA_TEMPR11[27] ), .Y(OR4_98_Y));
    OR4 OR4_321 (.A(\R_DATA_TEMPR0[5] ), .B(\R_DATA_TEMPR1[5] ), .C(
        \R_DATA_TEMPR2[5] ), .D(\R_DATA_TEMPR3[5] ), .Y(OR4_321_Y));
    OR4 OR4_615 (.A(\R_DATA_TEMPR8[75] ), .B(\R_DATA_TEMPR9[75] ), .C(
        \R_DATA_TEMPR10[75] ), .D(\R_DATA_TEMPR11[75] ), .Y(OR4_615_Y));
    OR4 OR4_337 (.A(\R_DATA_TEMPR8[71] ), .B(\R_DATA_TEMPR9[71] ), .C(
        \R_DATA_TEMPR10[71] ), .D(\R_DATA_TEMPR11[71] ), .Y(OR4_337_Y));
    OR4 OR4_130 (.A(\R_DATA_TEMPR16[35] ), .B(\R_DATA_TEMPR17[35] ), 
        .C(\R_DATA_TEMPR18[35] ), .D(\R_DATA_TEMPR19[35] ), .Y(
        OR4_130_Y));
    OR2 OR2_25 (.A(\R_DATA_TEMPR20[30] ), .B(\R_DATA_TEMPR21[30] ), .Y(
        OR2_25_Y));
    OR4 OR4_169 (.A(\R_DATA_TEMPR8[78] ), .B(\R_DATA_TEMPR9[78] ), .C(
        \R_DATA_TEMPR10[78] ), .D(\R_DATA_TEMPR11[78] ), .Y(OR4_169_Y));
    OR4 OR4_303 (.A(\R_DATA_TEMPR28[28] ), .B(\R_DATA_TEMPR29[28] ), 
        .C(\R_DATA_TEMPR30[28] ), .D(\R_DATA_TEMPR31[28] ), .Y(
        OR4_303_Y));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
