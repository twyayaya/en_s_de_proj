`timescale 1ns / 100ps


module error_gen(
    input [79:0] IN,
    output [79:0] OUT,
    input [63:0] selectt
    );
    
reg [79:0] IN_2;



always@(*) begin
    IN_2 = IN;
    case(selectt)
        64'd0  : IN_2[0] = ~IN[0] ;
        64'd1  : IN_2[1] = ~IN[1] ;
        64'd2  : IN_2[2] = ~IN[2] ;
        64'd3  : IN_2[3] = ~IN[3] ;
        64'd4  : IN_2[4] = ~IN[4] ;
        64'd5  : IN_2[5] = ~IN[5] ;
        64'd6  : IN_2[6] = ~IN[6] ;
        64'd7  : IN_2[7] = ~IN[7] ;
        64'd8  : IN_2[8] = ~IN[8] ;
        64'd9  : IN_2[9] = ~IN[9] ;
        64'd10  : IN_2[10] = ~IN[10] ;
        64'd11  : IN_2[11] = ~IN[11] ;
        64'd12  : IN_2[12] = ~IN[12] ;
        64'd13  : IN_2[13] = ~IN[13] ;
        64'd14  : IN_2[14] = ~IN[14] ;
        64'd15  : IN_2[15] = ~IN[15] ;
        64'd16  : IN_2[16] = ~IN[16] ;
        64'd17  : IN_2[17] = ~IN[17] ;
        64'd18  : IN_2[18] = ~IN[18] ;
        64'd19  : IN_2[19] = ~IN[19] ;
        64'd20  : IN_2[20] = ~IN[20] ;
        64'd21  : IN_2[21] = ~IN[21] ;
        64'd22  : IN_2[22] = ~IN[22] ;
        64'd23  : IN_2[23] = ~IN[23] ;
        64'd24  : IN_2[24] = ~IN[24] ;
        64'd25  : IN_2[25] = ~IN[25] ;
        64'd26  : IN_2[26] = ~IN[26] ;
        64'd27  : IN_2[27] = ~IN[27] ;
        64'd28  : IN_2[28] = ~IN[28] ;
        64'd29  : IN_2[29] = ~IN[29] ;
        64'd30  : IN_2[30] = ~IN[30] ;
        64'd31  : IN_2[31] = ~IN[31] ;
        64'd32  : IN_2[32] = ~IN[32] ;
        64'd33  : IN_2[33] = ~IN[33] ;
        64'd34  : IN_2[34] = ~IN[34] ;
        64'd35  : IN_2[35] = ~IN[35] ;
        64'd36  : IN_2[36] = ~IN[36] ;
        64'd37  : IN_2[37] = ~IN[37] ;
        64'd38  : IN_2[38] = ~IN[38] ;
        64'd39  : IN_2[39] = ~IN[39] ;
        64'd40  : IN_2[40] = ~IN[40] ;
        64'd41  : IN_2[41] = ~IN[41] ;
        64'd42  : IN_2[42] = ~IN[42] ;
        64'd43  : IN_2[43] = ~IN[43] ;
        64'd44  : IN_2[44] = ~IN[44] ;
        64'd45  : IN_2[45] = ~IN[45] ;
        64'd46  : IN_2[46] = ~IN[46] ;
        64'd47  : IN_2[47] = ~IN[47] ;
        64'd48  : IN_2[48] = ~IN[48] ;
        64'd49  : IN_2[49] = ~IN[49] ;
        64'd50  : IN_2[50] = ~IN[50] ;
        64'd51  : IN_2[51] = ~IN[51] ;
        64'd52  : IN_2[52] = ~IN[52] ;
        64'd53  : IN_2[53] = ~IN[53] ;
        64'd54  : IN_2[54] = ~IN[54] ;
        64'd55  : IN_2[55] = ~IN[55] ;
        64'd56  : IN_2[56] = ~IN[56] ;
        64'd57  : IN_2[57] = ~IN[57] ;
        64'd58  : IN_2[58] = ~IN[58] ;
        64'd59  : IN_2[59] = ~IN[59] ;
        64'd60  : IN_2[60] = ~IN[60] ;
        64'd61  : IN_2[61] = ~IN[61] ;
        64'd62  : IN_2[62] = ~IN[62] ;
        64'd63  : IN_2[63] = ~IN[63] ;
        
        default: IN_2 = IN ;
    endcase
end

assign OUT = IN_2;

endmodule