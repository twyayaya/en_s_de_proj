`timescale 1ns / 1ps

module de64_2 (
    input [71:0] INn, 
    input [7:0] SYNn,
    output [63:0] real_data

);

reg [71:0] LOC;
reg [71:0] OUT;
reg[63:0] r;

    always @(*) begin
        case(SYNn)
            8'b00100011: LOC <= 72'h00_0000_0000_0000_0001; 
            8'b01000011: LOC <= 72'h00_0000_0000_0000_0002;
            8'b10000011: LOC <= 72'h00_0000_0000_0000_0004;
            8'b00111101: LOC <= 72'h00_0000_0000_0000_0008;
            8'b01000101: LOC <= 72'h00_0000_0000_0000_0010;
            8'b10000101: LOC <= 72'h00_0000_0000_0000_0020;
            8'b10001001: LOC <= 72'h00_0000_0000_0000_0040;
            8'b01001001: LOC <= 72'h00_0000_0000_0000_0080;
            8'b01000110: LOC <= 72'h00_0000_0000_0000_0100;
            8'b10000110: LOC <= 72'h00_0000_0000_0000_0200;
            8'b00000111: LOC <= 72'h00_0000_0000_0000_0400;
            8'b01111010: LOC <= 72'h00_0000_0000_0000_0800;
            8'b10001010: LOC <= 72'h00_0000_0000_0000_1000;
            8'b00001011: LOC <= 72'h00_0000_0000_0000_2000;
            8'b00010011: LOC <= 72'h00_0000_0000_0000_4000;
            8'b10010010: LOC <= 72'h00_0000_0000_0000_8000;
            8'b10001100: LOC <= 72'h00_0000_0000_0001_0000;
            8'b00001101: LOC <= 72'h00_0000_0000_0002_0000;
            8'b00001110: LOC <= 72'h00_0000_0000_0004_0000;
            8'b11110100: LOC <= 72'h00_0000_0000_0008_0000;
            8'b00010101: LOC <= 72'h00_0000_0000_0010_0000;
            8'b00010110: LOC <= 72'h00_0000_0000_0020_0000;
            8'b00100110: LOC <= 72'h00_0000_0000_0040_0000;
            8'b00100101: LOC <= 72'h00_0000_0000_0080_0000;
            8'b00011001: LOC <= 72'h00_0000_0000_0100_0000;
            8'b00011010: LOC <= 72'h00_0000_0000_0200_0000;
            8'b00011100: LOC <= 72'h00_0000_0000_0400_0000;
            8'b11101001: LOC <= 72'h00_0000_0000_0800_0000;
            8'b00101010: LOC <= 72'h00_0000_0000_1000_0000;
            8'b00101100: LOC <= 72'h00_0000_0000_2000_0000;
            8'b01001100: LOC <= 72'h00_0000_0000_4000_0000;
            8'b01001010: LOC <= 72'h00_0000_0000_8000_0000;
            8'b00110010: LOC <= 72'h00_0000_0001_0000_0000;
            8'b00110100: LOC <= 72'h00_0000_0002_0000_0000;
            8'b00111000: LOC <= 72'h00_0000_0004_0000_0000;
            8'b11010011: LOC <= 72'h00_0000_0008_0000_0000;
            8'b01010100: LOC <= 72'h00_0000_0010_0000_0000;
            8'b01011000: LOC <= 72'h00_0000_0020_0000_0000;
            8'b10011000: LOC <= 72'h00_0000_0040_0000_0000;
            8'b10010100: LOC <= 72'h00_0000_0080_0000_0000;
            8'b01100100: LOC <= 72'h00_0000_0100_0000_0000;
            8'b01101000: LOC <= 72'h00_0000_0200_0000_0000;
            8'b01110000: LOC <= 72'h00_0000_0400_0000_0000;
            8'b10100111: LOC <= 72'h00_0000_0800_0000_0000;
            8'b10101000: LOC <= 72'h00_0000_1000_0000_0000;
            8'b10110000: LOC <= 72'h00_0000_2000_0000_0000;
            8'b00110001: LOC <= 72'h00_0000_4000_0000_0000;
            8'b00101001: LOC <= 72'h00_0000_8000_0000_0000;
            8'b11001000: LOC <= 72'h00_0001_0000_0000_0000;
            8'b11010000: LOC <= 72'h00_0002_0000_0000_0000;
            8'b11100000: LOC <= 72'h00_0004_0000_0000_0000;
            8'b01001111: LOC <= 72'h00_0008_0000_0000_0000;
            8'b01010001: LOC <= 72'h00_0010_0000_0000_0000;
            8'b01100001: LOC <= 72'h00_0020_0000_0000_0000;
            8'b01100010: LOC <= 72'h00_0040_0000_0000_0000;
            8'b01010010: LOC <= 72'h00_0080_0000_0000_0000;
            8'b10010001: LOC <= 72'h00_0100_0000_0000_0000;
            8'b10100001: LOC <= 72'h00_0200_0000_0000_0000;
            8'b11000001: LOC <= 72'h00_0400_0000_0000_0000;
            8'b10011110: LOC <= 72'h00_0800_0000_0000_0000;
            8'b10100010: LOC <= 72'h00_1000_0000_0000_0000;
            8'b11000010: LOC <= 72'h00_2000_0000_0000_0000;
            8'b11000100: LOC <= 72'h00_4000_0000_0000_0000;
            8'b10100100: LOC <= 72'h00_8000_0000_0000_0000;
            8'b00000001: LOC <= 72'h01_0000_0000_0000_0000;
            8'b00000010: LOC <= 72'h02_0000_0000_0000_0000;
            8'b00000100: LOC <= 72'h04_0000_0000_0000_0000;
            8'b00001000: LOC <= 72'h08_0000_0000_0000_0000;
            8'b00010000: LOC <= 72'h10_0000_0000_0000_0000;
            8'b00100000: LOC <= 72'h20_0000_0000_0000_0000;
            8'b01000000: LOC <= 72'h40_0000_0000_0000_0000;
            8'b10000000: LOC <= 72'h80_0000_0000_0000_0000;            
            default: LOC <= 0;
        endcase            
        OUT[71:0] <= LOC ^ INn[71:0];


        r = OUT[63:0];

    end
    

    assign real_data = r;
    

endmodule