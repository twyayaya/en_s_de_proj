`timescale 1 ns/100 ps
// Version: v12.5 12.900.11.2


module test6_for_compare(
       error_data_c,
       data_64_out_net_0,
       error_address_c,
       R_ADDR_c,
       ERRr_c
    );
output [63:0] error_data_c;
input  [63:0] data_64_out_net_0;
output [13:0] error_address_c;
input  [13:0] R_ADDR_c;
input  ERRr_c;

    wire GND, VCC;
    
    CFG2 #( .INIT(4'h8) )  \error_data[1]  (.A(ERRr_c), .B(
        data_64_out_net_0[1]), .Y(error_data_c[1]));
    CFG2 #( .INIT(4'h8) )  \error_data[43]  (.A(ERRr_c), .B(
        data_64_out_net_0[43]), .Y(error_data_c[43]));
    CFG2 #( .INIT(4'h8) )  \error_data[10]  (.A(ERRr_c), .B(
        data_64_out_net_0[10]), .Y(error_data_c[10]));
    CFG2 #( .INIT(4'h8) )  \error_data[50]  (.A(ERRr_c), .B(
        data_64_out_net_0[50]), .Y(error_data_c[50]));
    CFG2 #( .INIT(4'h8) )  \error_data[23]  (.A(ERRr_c), .B(
        data_64_out_net_0[23]), .Y(error_data_c[23]));
    CFG2 #( .INIT(4'h8) )  \error_data[36]  (.A(ERRr_c), .B(
        data_64_out_net_0[36]), .Y(error_data_c[36]));
    CFG2 #( .INIT(4'h8) )  \error_data[34]  (.A(ERRr_c), .B(
        data_64_out_net_0[34]), .Y(error_data_c[34]));
    CFG2 #( .INIT(4'h8) )  \error_data[37]  (.A(ERRr_c), .B(
        data_64_out_net_0[37]), .Y(error_data_c[37]));
    CFG2 #( .INIT(4'h8) )  \error_address[13]  (.A(ERRr_c), .B(
        R_ADDR_c[13]), .Y(error_address_c[13]));
    CFG2 #( .INIT(4'h8) )  \error_data[48]  (.A(ERRr_c), .B(
        data_64_out_net_0[48]), .Y(error_data_c[48]));
    CFG2 #( .INIT(4'h8) )  \error_address[12]  (.A(ERRr_c), .B(
        R_ADDR_c[12]), .Y(error_address_c[12]));
    CFG2 #( .INIT(4'h8) )  \error_data[49]  (.A(ERRr_c), .B(
        data_64_out_net_0[49]), .Y(error_data_c[49]));
    CFG2 #( .INIT(4'h8) )  \error_address[0]  (.A(ERRr_c), .B(
        R_ADDR_c[0]), .Y(error_address_c[0]));
    CFG2 #( .INIT(4'h8) )  \error_data[63]  (.A(ERRr_c), .B(
        data_64_out_net_0[63]), .Y(error_data_c[63]));
    CFG2 #( .INIT(4'h8) )  \error_data[2]  (.A(ERRr_c), .B(
        data_64_out_net_0[2]), .Y(error_data_c[2]));
    CFG2 #( .INIT(4'h8) )  \error_data[28]  (.A(ERRr_c), .B(
        data_64_out_net_0[28]), .Y(error_data_c[28]));
    CFG2 #( .INIT(4'h8) )  \error_data[45]  (.A(ERRr_c), .B(
        data_64_out_net_0[45]), .Y(error_data_c[45]));
    CFG2 #( .INIT(4'h8) )  \error_data[42]  (.A(ERRr_c), .B(
        data_64_out_net_0[42]), .Y(error_data_c[42]));
    CFG2 #( .INIT(4'h8) )  \error_address[11]  (.A(ERRr_c), .B(
        R_ADDR_c[11]), .Y(error_address_c[11]));
    CFG2 #( .INIT(4'h8) )  \error_data[41]  (.A(ERRr_c), .B(
        data_64_out_net_0[41]), .Y(error_data_c[41]));
    CFG2 #( .INIT(4'h8) )  \error_data[30]  (.A(ERRr_c), .B(
        data_64_out_net_0[30]), .Y(error_data_c[30]));
    CFG2 #( .INIT(4'h8) )  \error_data[29]  (.A(ERRr_c), .B(
        data_64_out_net_0[29]), .Y(error_data_c[29]));
    CFG2 #( .INIT(4'h8) )  \error_address[10]  (.A(ERRr_c), .B(
        R_ADDR_c[10]), .Y(error_address_c[10]));
    CFG2 #( .INIT(4'h8) )  \error_data[25]  (.A(ERRr_c), .B(
        data_64_out_net_0[25]), .Y(error_data_c[25]));
    CFG2 #( .INIT(4'h8) )  \error_data[22]  (.A(ERRr_c), .B(
        data_64_out_net_0[22]), .Y(error_data_c[22]));
    CFG2 #( .INIT(4'h8) )  \error_data[21]  (.A(ERRr_c), .B(
        data_64_out_net_0[21]), .Y(error_data_c[21]));
    CFG2 #( .INIT(4'h8) )  \error_data[3]  (.A(ERRr_c), .B(
        data_64_out_net_0[3]), .Y(error_data_c[3]));
    CFG2 #( .INIT(4'h8) )  \error_data[5]  (.A(ERRr_c), .B(
        data_64_out_net_0[5]), .Y(error_data_c[5]));
    CFG2 #( .INIT(4'h8) )  \error_address[9]  (.A(ERRr_c), .B(
        R_ADDR_c[9]), .Y(error_address_c[9]));
    CFG2 #( .INIT(4'h8) )  \error_data[46]  (.A(ERRr_c), .B(
        data_64_out_net_0[46]), .Y(error_data_c[46]));
    CFG2 #( .INIT(4'h8) )  \error_data[44]  (.A(ERRr_c), .B(
        data_64_out_net_0[44]), .Y(error_data_c[44]));
    CFG2 #( .INIT(4'h8) )  \error_data[7]  (.A(ERRr_c), .B(
        data_64_out_net_0[7]), .Y(error_data_c[7]));
    CFG2 #( .INIT(4'h8) )  \error_data[13]  (.A(ERRr_c), .B(
        data_64_out_net_0[13]), .Y(error_data_c[13]));
    CFG2 #( .INIT(4'h8) )  \error_data[53]  (.A(ERRr_c), .B(
        data_64_out_net_0[53]), .Y(error_data_c[53]));
    CFG2 #( .INIT(4'h8) )  \error_data[62]  (.A(ERRr_c), .B(
        data_64_out_net_0[62]), .Y(error_data_c[62]));
    CFG2 #( .INIT(4'h8) )  \error_data[47]  (.A(ERRr_c), .B(
        data_64_out_net_0[47]), .Y(error_data_c[47]));
    CFG2 #( .INIT(4'h8) )  \error_data[61]  (.A(ERRr_c), .B(
        data_64_out_net_0[61]), .Y(error_data_c[61]));
    CFG2 #( .INIT(4'h8) )  \error_data[26]  (.A(ERRr_c), .B(
        data_64_out_net_0[26]), .Y(error_data_c[26]));
    CFG2 #( .INIT(4'h8) )  \error_data[24]  (.A(ERRr_c), .B(
        data_64_out_net_0[24]), .Y(error_data_c[24]));
    CFG2 #( .INIT(4'h8) )  \error_data[27]  (.A(ERRr_c), .B(
        data_64_out_net_0[27]), .Y(error_data_c[27]));
    CFG2 #( .INIT(4'h8) )  \error_data[6]  (.A(ERRr_c), .B(
        data_64_out_net_0[6]), .Y(error_data_c[6]));
    CFG2 #( .INIT(4'h8) )  \error_address[4]  (.A(ERRr_c), .B(
        R_ADDR_c[4]), .Y(error_address_c[4]));
    CFG2 #( .INIT(4'h8) )  \error_address[8]  (.A(ERRr_c), .B(
        R_ADDR_c[8]), .Y(error_address_c[8]));
    CFG2 #( .INIT(4'h8) )  \error_address[2]  (.A(ERRr_c), .B(
        R_ADDR_c[2]), .Y(error_address_c[2]));
    CFG2 #( .INIT(4'h8) )  \error_data[8]  (.A(ERRr_c), .B(
        data_64_out_net_0[8]), .Y(error_data_c[8]));
    CFG2 #( .INIT(4'h8) )  \error_data[40]  (.A(ERRr_c), .B(
        data_64_out_net_0[40]), .Y(error_data_c[40]));
    CFG2 #( .INIT(4'h8) )  \error_data[9]  (.A(ERRr_c), .B(
        data_64_out_net_0[9]), .Y(error_data_c[9]));
    CFG2 #( .INIT(4'h8) )  \error_data[20]  (.A(ERRr_c), .B(
        data_64_out_net_0[20]), .Y(error_data_c[20]));
    CFG2 #( .INIT(4'h8) )  \error_data[4]  (.A(ERRr_c), .B(
        data_64_out_net_0[4]), .Y(error_data_c[4]));
    CFG2 #( .INIT(4'h8) )  \error_data[18]  (.A(ERRr_c), .B(
        data_64_out_net_0[18]), .Y(error_data_c[18]));
    GND GND_Z (.Y(GND));
    CFG2 #( .INIT(4'h8) )  \error_data[58]  (.A(ERRr_c), .B(
        data_64_out_net_0[58]), .Y(error_data_c[58]));
    VCC VCC_Z (.Y(VCC));
    CFG2 #( .INIT(4'h8) )  \error_data[19]  (.A(ERRr_c), .B(
        data_64_out_net_0[19]), .Y(error_data_c[19]));
    CFG2 #( .INIT(4'h8) )  \error_address[1]  (.A(ERRr_c), .B(
        R_ADDR_c[1]), .Y(error_address_c[1]));
    CFG2 #( .INIT(4'h8) )  \error_data[59]  (.A(ERRr_c), .B(
        data_64_out_net_0[59]), .Y(error_data_c[59]));
    CFG2 #( .INIT(4'h8) )  \error_data[33]  (.A(ERRr_c), .B(
        data_64_out_net_0[33]), .Y(error_data_c[33]));
    CFG2 #( .INIT(4'h8) )  \error_address[3]  (.A(ERRr_c), .B(
        R_ADDR_c[3]), .Y(error_address_c[3]));
    CFG2 #( .INIT(4'h8) )  \error_data[15]  (.A(ERRr_c), .B(
        data_64_out_net_0[15]), .Y(error_data_c[15]));
    CFG2 #( .INIT(4'h8) )  \error_data[12]  (.A(ERRr_c), .B(
        data_64_out_net_0[12]), .Y(error_data_c[12]));
    CFG2 #( .INIT(4'h8) )  \error_data[55]  (.A(ERRr_c), .B(
        data_64_out_net_0[55]), .Y(error_data_c[55]));
    CFG2 #( .INIT(4'h8) )  \error_data[52]  (.A(ERRr_c), .B(
        data_64_out_net_0[52]), .Y(error_data_c[52]));
    CFG2 #( .INIT(4'h8) )  \error_data[11]  (.A(ERRr_c), .B(
        data_64_out_net_0[11]), .Y(error_data_c[11]));
    CFG2 #( .INIT(4'h8) )  \error_data[51]  (.A(ERRr_c), .B(
        data_64_out_net_0[51]), .Y(error_data_c[51]));
    CFG2 #( .INIT(4'h8) )  \error_data[0]  (.A(ERRr_c), .B(
        data_64_out_net_0[0]), .Y(error_data_c[0]));
    CFG2 #( .INIT(4'h8) )  \error_address[7]  (.A(ERRr_c), .B(
        R_ADDR_c[7]), .Y(error_address_c[7]));
    CFG2 #( .INIT(4'h8) )  \error_data[60]  (.A(ERRr_c), .B(
        data_64_out_net_0[60]), .Y(error_data_c[60]));
    CFG2 #( .INIT(4'h8) )  \error_address[6]  (.A(ERRr_c), .B(
        R_ADDR_c[6]), .Y(error_address_c[6]));
    CFG2 #( .INIT(4'h8) )  \error_data[38]  (.A(ERRr_c), .B(
        data_64_out_net_0[38]), .Y(error_data_c[38]));
    CFG2 #( .INIT(4'h8) )  \error_data[39]  (.A(ERRr_c), .B(
        data_64_out_net_0[39]), .Y(error_data_c[39]));
    CFG2 #( .INIT(4'h8) )  \error_data[16]  (.A(ERRr_c), .B(
        data_64_out_net_0[16]), .Y(error_data_c[16]));
    CFG2 #( .INIT(4'h8) )  \error_data[14]  (.A(ERRr_c), .B(
        data_64_out_net_0[14]), .Y(error_data_c[14]));
    CFG2 #( .INIT(4'h8) )  \error_data[56]  (.A(ERRr_c), .B(
        data_64_out_net_0[56]), .Y(error_data_c[56]));
    CFG2 #( .INIT(4'h8) )  \error_data[54]  (.A(ERRr_c), .B(
        data_64_out_net_0[54]), .Y(error_data_c[54]));
    CFG2 #( .INIT(4'h8) )  \error_address[5]  (.A(ERRr_c), .B(
        R_ADDR_c[5]), .Y(error_address_c[5]));
    CFG2 #( .INIT(4'h8) )  \error_data[35]  (.A(ERRr_c), .B(
        data_64_out_net_0[35]), .Y(error_data_c[35]));
    CFG2 #( .INIT(4'h8) )  \error_data[32]  (.A(ERRr_c), .B(
        data_64_out_net_0[32]), .Y(error_data_c[32]));
    CFG2 #( .INIT(4'h8) )  \error_data[17]  (.A(ERRr_c), .B(
        data_64_out_net_0[17]), .Y(error_data_c[17]));
    CFG2 #( .INIT(4'h8) )  \error_data[57]  (.A(ERRr_c), .B(
        data_64_out_net_0[57]), .Y(error_data_c[57]));
    CFG2 #( .INIT(4'h8) )  \error_data[31]  (.A(ERRr_c), .B(
        data_64_out_net_0[31]), .Y(error_data_c[31]));
    
endmodule


module en64_RP2(
       en64_RP2_0_OUTt,
       W_DATA_c
    );
output [7:0] en64_RP2_0_OUTt;
input  [77:0] W_DATA_c;

    wire [5:5] OUTt_7_0_a2_6_a2_1;
    wire [0:0] OUTt_2_0_a2_0_a2_1_Z;
    wire [7:3] en64_RP2_0_OUTt_6;
    wire [1:1] OUTt_3_0_a2_0_a2_14_Z;
    wire [1:1] OUTt_3_0_a2_0_a2_10_Z;
    wire [1:1] OUTt_3_0_a2_0_a2_1_0_Z;
    wire [1:1] OUTt_3_0_a2_0_a2_4_Z;
    wire [5:5] OUTt_7_0_a2_6_a2_9_Z;
    wire [7:7] OUTt_1_0_a2_22_a2_9_Z;
    wire [7:7] OUTt_1_0_a2_22_a2_1;
    wire [0:0] OUTt_2_0_a2_0_a2_7_Z;
    wire [1:0] en64_RP2_0_OUTt_11;
    wire [3:3] en64_RP2_0_OUTt_3;
    wire [3:3] en64_RP2_0_OUTt_4;
    wire [3:3] en64_RP2_0_OUTt_5;
    wire [7:7] en64_RP2_0_OUTt_12;
    wire [6:6] OUTt_8_0_a2_13_Z;
    wire [6:6] OUTt_8_0_a2_12_Z;
    wire [6:6] OUTt_8_0_a2_11_Z;
    wire [6:6] OUTt_8_0_a2_1_Z;
    wire [6:6] OUTt_8_0_a2_0_Z;
    wire [0:0] OUTt_2_0_a2_0_a2_13_Z;
    wire [0:0] OUTt_2_0_a2_0_a2_12_Z;
    wire [0:0] OUTt_2_0_a2_0_a2_0_Z;
    wire [2:2] OUTt_4_0_a2_0_a2_11_Z;
    wire [2:2] OUTt_4_0_a2_0_a2_0_Z;
    wire [3:3] OUTt_5_0_a2_22_a2_12_Z;
    wire [3:3] OUTt_5_0_a2_22_a2_1_Z;
    wire [3:3] OUTt_5_0_a2_22_a2_0;
    wire [4:4] OUTt_6_0_a2_7_a2_14_Z;
    wire [4:4] OUTt_6_0_a2_7_a2_1;
    wire [4:4] OUTt_6_0_a2_7_a2_0;
    wire [5:5] OUTt_7_0_a2_6_a2_13_Z;
    wire [5:5] OUTt_7_0_a2_6_a2_12_Z;
    wire [5:5] OUTt_7_0_a2_6_a2_0_Z;
    wire [7:7] OUTt_1_0_a2_22_a2_13_Z;
    wire [7:7] OUTt_1_0_a2_22_a2_12_Z;
    wire [7:7] OUTt_1_0_a2_22_a2_0;
    wire [6:6] OUTt_8_0_a2_14_Z;
    wire [0:0] OUTt_2_0_a2_0_a2_14_Z;
    wire [1:1] OUTt_3_0_a2_0_a2_11_Z;
    wire [1:1] OUTt_3_0_a2_0_a2_8_Z;
    wire [2:2] OUTt_4_0_a2_0_a2_10_Z;
    wire [3:3] OUTt_5_0_a2_22_a2_11_Z;
    wire [3:3] OUTt_5_0_a2_22_a2_10_Z;
    wire [4:4] OUTt_6_0_a2_7_a2_13_Z;
    wire [4:4] OUTt_6_0_a2_7_a2_12_Z;
    wire [5:5] OUTt_7_0_a2_6_a2_14_Z;
    wire [7:7] OUTt_1_0_a2_22_a2_14_Z;
    wire [6:6] OUTt_8_0_a2_15_Z;
    wire [0:0] OUTt_2_0_a2_0_a2_16_Z;
    wire [0:0] OUTt_2_0_a2_0_a2_15_Z;
    wire [2:2] OUTt_4_0_a2_0_a2_12_Z;
    wire [3:3] OUTt_5_0_a2_22_a2_13_Z;
    wire [4:4] OUTt_6_0_a2_7_a2_16_Z;
    wire [4:4] OUTt_6_0_a2_7_a2_15_Z;
    wire [5:5] OUTt_7_0_a2_6_a2_18_Z;
    wire [5:5] OUTt_7_0_a2_6_a2_16_Z;
    wire [7:7] OUTt_1_0_a2_22_a2_18_Z;
    wire [7:7] OUTt_1_0_a2_22_a2_16_Z;
    wire [2:2] OUTt_4_0_a2_0_a2_9_Z;
    wire N_3, GND, VCC;
    
    CFG4 #( .INIT(16'h6996) )  \OUTt_5_0_a2_22_a2_10[3]  (.A(
        en64_RP2_0_OUTt_4[3]), .B(en64_RP2_0_OUTt_3[3]), .C(
        W_DATA_c[37]), .D(W_DATA_c[35]), .Y(OUTt_5_0_a2_22_a2_10_Z[3]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_5_0_a2_22_a2_12[3]  (.A(
        W_DATA_c[57]), .B(W_DATA_c[51]), .C(W_DATA_c[46]), .D(
        W_DATA_c[42]), .Y(OUTt_5_0_a2_22_a2_12_Z[3]));
    CFG2 #( .INIT(4'h6) )  \OUTt_5_0_a2_22_a2_5[3]  (.A(W_DATA_c[20]), 
        .B(W_DATA_c[21]), .Y(en64_RP2_0_OUTt_5[3]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_2_0_a2_0_a2_13[0]  (.A(
        W_DATA_c[72]), .B(W_DATA_c[16]), .C(W_DATA_c[15]), .D(
        W_DATA_c[12]), .Y(OUTt_2_0_a2_0_a2_13_Z[0]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_1_0_a2_22_a2_14[7]  (.A(
        en64_RP2_0_OUTt_12[7]), .B(en64_RP2_0_OUTt_6[7]), .C(
        W_DATA_c[23]), .D(W_DATA_c[20]), .Y(OUTt_1_0_a2_22_a2_14_Z[7]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_7_0_a2_6_a2_16[5]  (.A(
        OUTt_7_0_a2_6_a2_1[5]), .B(OUTt_7_0_a2_6_a2_0_Z[5]), .C(
        W_DATA_c[62]), .D(W_DATA_c[57]), .Y(OUTt_7_0_a2_6_a2_16_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_6_0_a2_7_a2_14[4]  (.A(
        W_DATA_c[70]), .B(W_DATA_c[67]), .C(W_DATA_c[64]), .D(
        W_DATA_c[56]), .Y(OUTt_6_0_a2_7_a2_14_Z[4]));
    CFG2 #( .INIT(4'h6) )  \OUTt_2_0_a2_0_a2_11[0]  (.A(W_DATA_c[64]), 
        .B(W_DATA_c[65]), .Y(en64_RP2_0_OUTt_11[0]));
    CFG3 #( .INIT(8'h96) )  \OUTt_7_0_a2_6_a2_0_0[5]  (.A(W_DATA_c[50])
        , .B(W_DATA_c[23]), .C(W_DATA_c[0]), .Y(
        OUTt_7_0_a2_6_a2_0_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_2_0_a2_0_a2_12[0]  (.A(
        W_DATA_c[43]), .B(W_DATA_c[27]), .C(W_DATA_c[24]), .D(
        W_DATA_c[21]), .Y(OUTt_2_0_a2_0_a2_12_Z[0]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_8_0_a2_0[6]  (.A(W_DATA_c[75]), 
        .B(W_DATA_c[63]), .C(W_DATA_c[43]), .D(W_DATA_c[36]), .Y(
        OUTt_8_0_a2_0_Z[6]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_5_0_a2_22_a2_11[3]  (.A(
        en64_RP2_0_OUTt_6[3]), .B(en64_RP2_0_OUTt_5[3]), .C(
        W_DATA_c[34]), .D(W_DATA_c[32]), .Y(OUTt_5_0_a2_22_a2_11_Z[3]));
    CFG2 #( .INIT(4'h6) )  \OUTt_5_0_a2_22_a2_6[3]  (.A(W_DATA_c[22]), 
        .B(W_DATA_c[31]), .Y(en64_RP2_0_OUTt_6[3]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_7_0_a2_6_a2[5]  (.A(
        OUTt_7_0_a2_6_a2_18_Z[5]), .B(OUTt_7_0_a2_6_a2_16_Z[5]), .C(
        OUTt_7_0_a2_6_a2_13_Z[5]), .D(OUTt_7_0_a2_6_a2_12_Z[5]), .Y(
        en64_RP2_0_OUTt[5]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_4_0_a2_0_a2_12[2]  (.A(
        en64_RP2_0_OUTt_12[7]), .B(OUTt_4_0_a2_0_a2_0_Z[2]), .C(
        W_DATA_c[41]), .D(W_DATA_c[35]), .Y(OUTt_4_0_a2_0_a2_12_Z[2]));
    CFG2 #( .INIT(4'h6) )  \OUTt_1_0_a2_22_a2_12[7]  (.A(W_DATA_c[76]), 
        .B(W_DATA_c[77]), .Y(en64_RP2_0_OUTt_12[7]));
    CFG2 #( .INIT(4'h6) )  \OUTt_1_0_a2_22_a2_6[7]  (.A(W_DATA_c[46]), 
        .B(W_DATA_c[47]), .Y(en64_RP2_0_OUTt_6[7]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_8_0_a2[6]  (.A(
        OUTt_8_0_a2_15_Z[6]), .B(OUTt_8_0_a2_14_Z[6]), .C(
        OUTt_8_0_a2_13_Z[6]), .D(OUTt_8_0_a2_12_Z[6]), .Y(
        en64_RP2_0_OUTt[6]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_4_0_a2_0_a2_9[2]  (.A(
        OUTt_3_0_a2_0_a2_4_Z[1]), .B(OUTt_2_0_a2_0_a2_7_Z[0]), .C(
        W_DATA_c[32]), .D(W_DATA_c[3]), .Y(OUTt_4_0_a2_0_a2_9_Z[2]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_3_0_a2_0_a2[1]  (.A(
        en64_RP2_0_OUTt_6[3]), .B(OUTt_3_0_a2_0_a2_14_Z[1]), .C(
        OUTt_3_0_a2_0_a2_10_Z[1]), .D(OUTt_3_0_a2_0_a2_1_0_Z[1]), .Y(
        en64_RP2_0_OUTt[1]));
    CFG2 #( .INIT(4'h6) )  \OUTt_2_0_a2_0_a2_7[0]  (.A(W_DATA_c[4]), 
        .B(W_DATA_c[5]), .Y(OUTt_2_0_a2_0_a2_7_Z[0]));
    CFG3 #( .INIT(8'h96) )  \OUTt_2_0_a2_0_a2_0[0]  (.A(W_DATA_c[30]), 
        .B(W_DATA_c[3]), .C(W_DATA_c[0]), .Y(OUTt_2_0_a2_0_a2_0_Z[0]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_6_0_a2_7_a2_13[4]  (.A(
        en64_RP2_0_OUTt_6[5]), .B(W_DATA_c[43]), .C(W_DATA_c[40]), .D(
        W_DATA_c[32]), .Y(OUTt_6_0_a2_7_a2_13_Z[4]));
    CFG2 #( .INIT(4'h6) )  \OUTt_5_0_a2_22_a2_3[3]  (.A(W_DATA_c[6]), 
        .B(W_DATA_c[7]), .Y(en64_RP2_0_OUTt_3[3]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_2_0_a2_0_a2_1[0]  (.A(W_DATA_c[6])
        , .B(W_DATA_c[7]), .C(W_DATA_c[1]), .D(W_DATA_c[2]), .Y(
        OUTt_2_0_a2_0_a2_1_Z[0]));
    CFG2 #( .INIT(4'h6) )  \OUTt_5_0_a2_22_a2_4[3]  (.A(W_DATA_c[14]), 
        .B(W_DATA_c[15]), .Y(en64_RP2_0_OUTt_4[3]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_6_0_a2_7_a2_1_0[4]  (.A(
        W_DATA_c[73]), .B(W_DATA_c[45]), .C(W_DATA_c[25]), .D(
        W_DATA_c[13]), .Y(OUTt_6_0_a2_7_a2_1[4]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_3_0_a2_0_a2_11_0[1]  (.A(
        en64_RP2_0_OUTt_11[1]), .B(W_DATA_c[74]), .C(W_DATA_c[63]), .D(
        W_DATA_c[13]), .Y(OUTt_3_0_a2_0_a2_11_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_8_0_a2_14[6]  (.A(
        en64_RP2_0_OUTt_11[1]), .B(en64_RP2_0_OUTt_11[0]), .C(
        W_DATA_c[76]), .D(W_DATA_c[72]), .Y(OUTt_8_0_a2_14_Z[6]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_1_0_a2_22_a2_13[7]  (.A(
        W_DATA_c[61]), .B(W_DATA_c[60]), .C(W_DATA_c[55]), .D(
        W_DATA_c[53]), .Y(OUTt_1_0_a2_22_a2_13_Z[7]));
    CFG3 #( .INIT(8'h96) )  \OUTt_8_0_a2_15[6]  (.A(
        OUTt_8_0_a2_11_Z[6]), .B(OUTt_8_0_a2_1_Z[6]), .C(
        OUTt_8_0_a2_0_Z[6]), .Y(OUTt_8_0_a2_15_Z[6]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_4_0_a2_0_a2_10[2]  (.A(
        en64_RP2_0_OUTt_5[3]), .B(W_DATA_c[27]), .C(W_DATA_c[24]), .D(
        W_DATA_c[22]), .Y(OUTt_4_0_a2_0_a2_10_Z[2]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_3_0_a2_0_a2_8[1]  (.A(
        W_DATA_c[75]), .B(W_DATA_c[43]), .C(W_DATA_c[34]), .D(
        W_DATA_c[0]), .Y(OUTt_3_0_a2_0_a2_8_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_2_0_a2_0_a2[0]  (.A(
        OUTt_2_0_a2_0_a2_16_Z[0]), .B(OUTt_2_0_a2_0_a2_15_Z[0]), .C(
        OUTt_2_0_a2_0_a2_14_Z[0]), .D(OUTt_2_0_a2_0_a2_13_Z[0]), .Y(
        en64_RP2_0_OUTt[0]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_8_0_a2_12[6]  (.A(W_DATA_c[62]), 
        .B(W_DATA_c[61]), .C(W_DATA_c[60]), .D(W_DATA_c[52]), .Y(
        OUTt_8_0_a2_12_Z[6]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_7_0_a2_6_a2_14[5]  (.A(
        en64_RP2_0_OUTt_6[5]), .B(W_DATA_c[77]), .C(W_DATA_c[40]), .D(
        W_DATA_c[35]), .Y(OUTt_7_0_a2_6_a2_14_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_5_0_a2_22_a2_1[3]  (.A(
        W_DATA_c[54]), .B(W_DATA_c[45]), .C(W_DATA_c[33]), .D(
        W_DATA_c[13]), .Y(OUTt_5_0_a2_22_a2_1_Z[3]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_6_0_a2_7_a2_15[4]  (.A(
        OUTt_6_0_a2_7_a2_0[4]), .B(W_DATA_c[61]), .C(W_DATA_c[55]), .D(
        W_DATA_c[52]), .Y(OUTt_6_0_a2_7_a2_15_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_5_0_a2_22_a2[3]  (.A(
        OUTt_5_0_a2_22_a2_13_Z[3]), .B(OUTt_5_0_a2_22_a2_12_Z[3]), .C(
        OUTt_5_0_a2_22_a2_11_Z[3]), .D(OUTt_5_0_a2_22_a2_10_Z[3]), .Y(
        en64_RP2_0_OUTt[3]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_2_0_a2_0_a2_16[0]  (.A(
        OUTt_2_0_a2_0_a2_12_Z[0]), .B(OUTt_2_0_a2_0_a2_7_Z[0]), .C(
        OUTt_2_0_a2_0_a2_1_Z[0]), .D(W_DATA_c[33]), .Y(
        OUTt_2_0_a2_0_a2_16_Z[0]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_2_0_a2_0_a2_14[0]  (.A(
        en64_RP2_0_OUTt_11[0]), .B(W_DATA_c[71]), .C(W_DATA_c[70]), .D(
        W_DATA_c[63]), .Y(OUTt_2_0_a2_0_a2_14_Z[0]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_1_0_a2_22_a2_16[7]  (.A(
        OUTt_1_0_a2_22_a2_1[7]), .B(OUTt_1_0_a2_22_a2_0[7]), .C(
        W_DATA_c[70]), .D(W_DATA_c[62]), .Y(OUTt_1_0_a2_22_a2_16_Z[7]));
    CFG2 #( .INIT(4'h6) )  \OUTt_1_0_a2_22_a2_9[7]  (.A(W_DATA_c[71]), 
        .B(W_DATA_c[72]), .Y(OUTt_1_0_a2_22_a2_9_Z[7]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_2_0_a2_0_a2_15[0]  (.A(
        OUTt_2_0_a2_0_a2_0_Z[0]), .B(W_DATA_c[57]), .C(W_DATA_c[56]), 
        .D(W_DATA_c[53]), .Y(OUTt_2_0_a2_0_a2_15_Z[0]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_3_0_a2_0_a2_10[1]  (.A(
        en64_RP2_0_OUTt_4[3]), .B(W_DATA_c[17]), .C(W_DATA_c[16]), .D(
        W_DATA_c[12]), .Y(OUTt_3_0_a2_0_a2_10_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_8_0_a2_11[6]  (.A(W_DATA_c[10]), 
        .B(W_DATA_c[7]), .C(W_DATA_c[4]), .D(W_DATA_c[1]), .Y(
        OUTt_8_0_a2_11_Z[6]));
    CFG2 #( .INIT(4'h6) )  \OUTt_7_0_a2_6_a2_6[5]  (.A(W_DATA_c[41]), 
        .B(W_DATA_c[42]), .Y(en64_RP2_0_OUTt_6[5]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_7_0_a2_6_a2_12[5]  (.A(
        W_DATA_c[34]), .B(W_DATA_c[27]), .C(W_DATA_c[13]), .D(
        W_DATA_c[3]), .Y(OUTt_7_0_a2_6_a2_12_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_5_0_a2_22_a2_0_0[3]  (.A(
        W_DATA_c[63]), .B(W_DATA_c[36]), .C(W_DATA_c[30]), .D(
        W_DATA_c[3]), .Y(OUTt_5_0_a2_22_a2_0[3]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_3_0_a2_0_a2_4[1]  (.A(
        W_DATA_c[73]), .B(W_DATA_c[25]), .C(W_DATA_c[10]), .D(N_3), .Y(
        OUTt_3_0_a2_0_a2_4_Z[1]));
    CFG2 #( .INIT(4'h6) )  \OUTt_1_0_a2_22_a2_1_0[7]  (.A(W_DATA_c[2]), 
        .B(W_DATA_c[5]), .Y(OUTt_1_0_a2_22_a2_1[7]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_8_0_a2_1[6]  (.A(W_DATA_c[50]), 
        .B(W_DATA_c[45]), .C(W_DATA_c[23]), .D(W_DATA_c[13]), .Y(
        OUTt_8_0_a2_1_Z[6]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_5_0_a2_22_a2_13[3]  (.A(
        OUTt_5_0_a2_22_a2_1_Z[3]), .B(OUTt_5_0_a2_22_a2_0[3]), .C(
        W_DATA_c[73]), .D(W_DATA_c[60]), .Y(OUTt_5_0_a2_22_a2_13_Z[3]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_7_0_a2_6_a2_18[5]  (.A(
        OUTt_7_0_a2_6_a2_14_Z[5]), .B(OUTt_7_0_a2_6_a2_9_Z[5]), .C(
        W_DATA_c[74]), .D(W_DATA_c[71]), .Y(OUTt_7_0_a2_6_a2_18_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_6_0_a2_7_a2_12[4]  (.A(
        en64_RP2_0_OUTt_6[7]), .B(W_DATA_c[44]), .C(W_DATA_c[23]), .D(
        W_DATA_c[17]), .Y(OUTt_6_0_a2_7_a2_12_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_4_0_a2_0_a2_11[2]  (.A(
        W_DATA_c[47]), .B(W_DATA_c[44]), .C(W_DATA_c[12]), .D(
        W_DATA_c[11]), .Y(OUTt_4_0_a2_0_a2_11_Z[2]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_1_0_a2_22_a2[7]  (.A(
        OUTt_1_0_a2_22_a2_18_Z[7]), .B(OUTt_1_0_a2_22_a2_16_Z[7]), .C(
        OUTt_1_0_a2_22_a2_13_Z[7]), .D(OUTt_1_0_a2_22_a2_12_Z[7]), .Y(
        en64_RP2_0_OUTt[7]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_6_0_a2_7_a2_16[4]  (.A(
        OUTt_6_0_a2_7_a2_12_Z[4]), .B(OUTt_6_0_a2_7_a2_1[4]), .C(
        W_DATA_c[31]), .D(W_DATA_c[24]), .Y(OUTt_6_0_a2_7_a2_16_Z[4]));
    GND GND_Z (.Y(GND));
    VCC VCC_Z (.Y(VCC));
    CFG2 #( .INIT(4'h6) )  \OUTt_3_0_a2_0_a2_11[1]  (.A(W_DATA_c[66]), 
        .B(W_DATA_c[67]), .Y(en64_RP2_0_OUTt_11[1]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_1_0_a2_22_a2_0_0[7]  (.A(
        W_DATA_c[75]), .B(W_DATA_c[54]), .C(W_DATA_c[43]), .D(
        W_DATA_c[33]), .Y(OUTt_1_0_a2_22_a2_0[7]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_3_0_a2_0_a2_1_0[1]  (.A(
        OUTt_3_0_a2_0_a2_4_Z[1]), .B(W_DATA_c[11]), .C(W_DATA_c[2]), 
        .D(W_DATA_c[1]), .Y(OUTt_3_0_a2_0_a2_1_0_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_8_0_a2_13[6]  (.A(W_DATA_c[51]), 
        .B(W_DATA_c[44]), .C(W_DATA_c[37]), .D(W_DATA_c[33]), .Y(
        OUTt_8_0_a2_13_Z[6]));
    CFG3 #( .INIT(8'h96) )  \OUTt_6_0_a2_7_a2_0_0[4]  (.A(W_DATA_c[30])
        , .B(W_DATA_c[16]), .C(W_DATA_c[3]), .Y(OUTt_6_0_a2_7_a2_0[4]));
    CFG2 #( .INIT(4'h6) )  \OUTt_7_0_a2_6_a2_9[5]  (.A(W_DATA_c[65]), 
        .B(W_DATA_c[66]), .Y(OUTt_7_0_a2_6_a2_9_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_7_0_a2_6_a2_13[5]  (.A(
        W_DATA_c[56]), .B(W_DATA_c[55]), .C(W_DATA_c[52]), .D(
        W_DATA_c[51]), .Y(OUTt_7_0_a2_6_a2_13_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_4_0_a2_0_a2[2]  (.A(
        OUTt_4_0_a2_0_a2_12_Z[2]), .B(OUTt_4_0_a2_0_a2_11_Z[2]), .C(
        OUTt_4_0_a2_0_a2_10_Z[2]), .D(OUTt_4_0_a2_0_a2_9_Z[2]), .Y(
        en64_RP2_0_OUTt[2]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_1_0_a2_22_a2_12_0[7]  (.A(
        W_DATA_c[17]), .B(W_DATA_c[14]), .C(W_DATA_c[11]), .D(
        W_DATA_c[6]), .Y(OUTt_1_0_a2_22_a2_12_Z[7]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_1_0_a2_22_a2_18[7]  (.A(
        OUTt_1_0_a2_22_a2_14_Z[7]), .B(OUTt_1_0_a2_22_a2_9_Z[7]), .C(
        W_DATA_c[74]), .D(W_DATA_c[73]), .Y(OUTt_1_0_a2_22_a2_18_Z[7]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_3_0_a2_0_a2_14[1]  (.A(
        OUTt_3_0_a2_0_a2_11_Z[1]), .B(OUTt_3_0_a2_0_a2_8_Z[1]), .C(
        W_DATA_c[40]), .D(W_DATA_c[37]), .Y(OUTt_3_0_a2_0_a2_14_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_7_0_a2_6_a2_1_0[5]  (.A(
        W_DATA_c[26]), .B(W_DATA_c[53]), .C(W_DATA_c[33]), .D(
        W_DATA_c[54]), .Y(OUTt_7_0_a2_6_a2_1[5]));
    CFG2 #( .INIT(4'h6) )  \OUTt_7_0_a2_6_a2_0[5]  (.A(W_DATA_c[26]), 
        .B(W_DATA_c[53]), .Y(N_3));
    CFG4 #( .INIT(16'h6996) )  \OUTt_6_0_a2_7_a2[4]  (.A(
        OUTt_6_0_a2_7_a2_16_Z[4]), .B(OUTt_6_0_a2_7_a2_15_Z[4]), .C(
        OUTt_6_0_a2_7_a2_14_Z[4]), .D(OUTt_6_0_a2_7_a2_13_Z[4]), .Y(
        en64_RP2_0_OUTt[4]));
    CFG4 #( .INIT(16'h6996) )  \OUTt_4_0_a2_0_a2_0[2]  (.A(
        W_DATA_c[63]), .B(W_DATA_c[50]), .C(W_DATA_c[36]), .D(
        W_DATA_c[23]), .Y(OUTt_4_0_a2_0_a2_0_Z[2]));
    
endmodule


module de64_1(
       PF_TPSRAM_C0_0_R_DATA,
       data_64_out_net_0,
       ERRr_c
    );
input  [7:0] PF_TPSRAM_C0_0_R_DATA;
input  [63:0] data_64_out_net_0;
output ERRr_c;

    wire [3:3] SYN_5_0_a2_7_Z;
    wire [4:4] SYN_6_0_Z;
    wire [7:7] SYN_1;
    wire [1:1] SYN_3_0_a2_0_Z;
    wire [0:0] SYN_2_0_a2_0_Z;
    wire [2:2] SYN_4_0_a2_10_Z;
    wire [2:2] SYN_4_0_a2_15_Z;
    wire [4:4] SYN_6_8_Z;
    wire [2:2] SYN_4_0_a2_1_Z;
    wire [5:5] SYN_7_0_a2_6_Z;
    wire [1:1] SYN_3_0_a2_4_Z;
    wire [4:4] SYN_6_3_0;
    wire [4:4] SYN_6_12_Z;
    wire [7:7] SYN_6;
    wire [7:6] SYN_8;
    wire [4:4] SYN_6_3_Z;
    wire [2:2] SYN_4_5;
    wire [1:1] SYN_3_5;
    wire [4:4] SYN_6_12_0_Z;
    wire [4:4] SYN_6_11_Z;
    wire [0:0] SYN_2_0_a2_13_Z;
    wire [0:0] SYN_2_0_a2_12_Z;
    wire [0:0] SYN_2_0_a2_11_Z;
    wire [0:0] SYN_2_0_a2_9;
    wire [1:1] SYN_3_0_a2_12_Z;
    wire [1:1] SYN_3_0_a2_10_Z;
    wire [2:2] SYN_4_0_a2_14_Z;
    wire [2:2] SYN_4_0_a2_12_Z;
    wire [3:3] SYN_5_0_a2_12_Z;
    wire [3:3] SYN_5_0_a2_11_Z;
    wire [5:5] SYN_7_0_a2_14_Z;
    wire [5:5] SYN_7_0_a2_12_Z;
    wire [5:5] SYN_7_0_a2_2_Z;
    wire [6:6] SYN_8_0_a2_10_Z;
    wire [6:6] SYN_8_0_a2_1;
    wire [7:7] SYN_0_a2_12_Z;
    wire [7:7] SYN_0_a2_3_Z;
    wire [0:0] SYN_2_14;
    wire [4:4] SYN_6_4_Z;
    wire [1:1] SYN_3_10;
    wire [1:1] SYN_3_0_a2_15_Z;
    wire [2:2] SYN_4_0_a2_13_Z;
    wire [3:3] SYN_5_0_a2_10_Z;
    wire [5:5] SYN_7_0_a2_11_Z;
    wire [5:5] SYN_7_0_a2_10_Z;
    wire [6:6] SYN_8_0_a2_12_Z;
    wire [6:6] SYN_8_0_a2_11_Z;
    wire [6:6] SYN_8_0_a2_9_Z;
    wire [7:7] SYN_0_a2_13_Z;
    wire [7:7] SYN_0_a2_10_Z;
    wire [4:4] SYN_6_15_Z;
    wire [4:4] SYN_6_13_Z;
    wire [0:0] SYN_2_0_a2_15_Z;
    wire [0:0] SYN_2_0_a2_14_Z;
    wire [1:1] SYN_3_0_a2_13_Z;
    wire [2:2] SYN_4_0_a2_16_Z;
    wire [3:3] SYN_5_0_a2_16_Z;
    wire [3:3] SYN_5_0_a2_14_Z;
    wire [6:6] SYN_8_0_a2_13_Z;
    wire [7:7] SYN_0_a2_15_Z;
    wire [7:7] SYN_0_a2_9_Z;
    wire [4:4] SYN_6_17_Z;
    wire [5:5] SYN_7_0_a2_16_Z;
    wire [1:1] SYN_3_0_a2_16_Z;
    wire [5:5] SYN_7;
    wire [3:3] SYN_5;
    wire [2:2] SYN_4;
    wire [0:0] SYN_2;
    wire [4:4] SYN_6_Z;
    wire [7:7] SYN;
    wire N_31, N_32, N_27, ERRr_4_Z, ERRr_2_Z, GND, VCC;
    
    CFG4 #( .INIT(16'h6996) )  \SYN_4_0_a2[2]  (.A(SYN_4_0_a2_16_Z[2]), 
        .B(SYN_4_0_a2_15_Z[2]), .C(SYN_4_0_a2_14_Z[2]), .D(
        SYN_4_0_a2_13_Z[2]), .Y(SYN_4[2]));
    CFG4 #( .INIT(16'h6996) )  \SYN_2_0_a2_15[0]  (.A(
        SYN_2_0_a2_11_Z[0]), .B(SYN_2_0_a2_0_Z[0]), .C(
        data_64_out_net_0[2]), .D(PF_TPSRAM_C0_0_R_DATA[0]), .Y(
        SYN_2_0_a2_15_Z[0]));
    CFG3 #( .INIT(8'h96) )  \SYN_2_0_a2_14_0[0]  (.A(SYN_2_14[0]), .B(
        SYN_2_0_a2_9[0]), .C(data_64_out_net_0[58]), .Y(
        SYN_2_0_a2_14_Z[0]));
    CFG2 #( .INIT(4'h6) )  \SYN_5_0_a2_1[3]  (.A(data_64_out_net_0[25])
        , .B(data_64_out_net_0[26]), .Y(SYN_6_3_0[4]));
    CFG2 #( .INIT(4'h6) )  \SYN_0_a2_1[7]  (.A(data_64_out_net_0[12]), 
        .B(data_64_out_net_0[59]), .Y(N_31));
    CFG4 #( .INIT(16'h6996) )  \SYN_2_0_a2[0]  (.A(SYN_2_0_a2_15_Z[0]), 
        .B(SYN_2_0_a2_14_Z[0]), .C(SYN_2_0_a2_13_Z[0]), .D(
        SYN_2_0_a2_12_Z[0]), .Y(SYN_2[0]));
    CFG2 #( .INIT(4'h6) )  \SYN_6_3[4]  (.A(data_64_out_net_0[15]), .B(
        data_64_out_net_0[19]), .Y(SYN_6_3_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \SYN_7_0_a2_10[5]  (.A(
        data_64_out_net_0[23]), .B(data_64_out_net_0[22]), .C(
        PF_TPSRAM_C0_0_R_DATA[5]), .D(N_32), .Y(SYN_7_0_a2_10_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \SYN_5_0_a2_12[3]  (.A(
        data_64_out_net_0[37]), .B(data_64_out_net_0[34]), .C(
        data_64_out_net_0[31]), .D(data_64_out_net_0[30]), .Y(
        SYN_5_0_a2_12_Z[3]));
    CFG4 #( .INIT(16'h6996) )  \SYN_4_0_a2_10[2]  (.A(SYN_3_5[1]), .B(
        data_64_out_net_0[51]), .C(data_64_out_net_0[8]), .D(
        PF_TPSRAM_C0_0_R_DATA[2]), .Y(SYN_4_0_a2_10_Z[2]));
    CFG4 #( .INIT(16'hFFFE) )  ERRr_4 (.A(SYN_8[6]), .B(SYN_7[5]), .C(
        SYN_6_Z[4]), .D(SYN_4[2]), .Y(ERRr_4_Z));
    CFG3 #( .INIT(8'hBE) )  ERRr_2 (.A(SYN_5[3]), .B(
        SYN_3_0_a2_16_Z[1]), .C(SYN_3_0_a2_15_Z[1]), .Y(ERRr_2_Z));
    CFG4 #( .INIT(16'h6996) )  \SYN_6_12_0[4]  (.A(
        data_64_out_net_0[59]), .B(data_64_out_net_0[56]), .C(
        data_64_out_net_0[55]), .D(data_64_out_net_0[38]), .Y(
        SYN_6_12_0_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \SYN_7_0_a2_16[5]  (.A(
        SYN_7_0_a2_12_Z[5]), .B(SYN_7_0_a2_6_Z[5]), .C(
        data_64_out_net_0[57]), .D(data_64_out_net_0[50]), .Y(
        SYN_7_0_a2_16_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \SYN_3_0_a2_13[1]  (.A(SYN_3_10[1]), .B(
        SYN_3_5[1]), .C(data_64_out_net_0[55]), .D(
        data_64_out_net_0[13]), .Y(SYN_3_0_a2_13_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \SYN_6[4]  (.A(SYN_6_17_Z[4]), .B(
        SYN_6_15_Z[4]), .C(SYN_6_12_0_Z[4]), .D(SYN_6_11_Z[4]), .Y(
        SYN_6_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \SYN_3_0_a2_10_0[1]  (.A(
        data_64_out_net_0[10]), .B(data_64_out_net_0[9]), .C(
        data_64_out_net_0[2]), .D(PF_TPSRAM_C0_0_R_DATA[1]), .Y(
        SYN_3_0_a2_10_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \SYN_8_0_a2[6]  (.A(SYN_8_0_a2_13_Z[6]), 
        .B(SYN_8_0_a2_12_Z[6]), .C(SYN_8_0_a2_11_Z[6]), .D(
        SYN_8_0_a2_10_Z[6]), .Y(SYN_8[6]));
    CFG4 #( .INIT(16'h6996) )  \SYN_0_a2_9[7]  (.A(SYN_1[7]), .B(
        data_64_out_net_0[48]), .C(data_64_out_net_0[44]), .D(
        data_64_out_net_0[2]), .Y(SYN_0_a2_9_Z[7]));
    CFG4 #( .INIT(16'h6996) )  \SYN_8_0_a2_12[6]  (.A(SYN_6[7]), .B(
        data_64_out_net_0[48]), .C(data_64_out_net_0[41]), .D(
        data_64_out_net_0[37]), .Y(SYN_8_0_a2_12_Z[6]));
    CFG4 #( .INIT(16'h6996) )  \SYN_5_0_a2_11[3]  (.A(
        data_64_out_net_0[18]), .B(data_64_out_net_0[17]), .C(
        data_64_out_net_0[16]), .D(data_64_out_net_0[13]), .Y(
        SYN_5_0_a2_11_Z[3]));
    CFG4 #( .INIT(16'h6996) )  \SYN_3_0_a2_12[1]  (.A(
        data_64_out_net_0[28]), .B(data_64_out_net_0[21]), .C(
        data_64_out_net_0[15]), .D(data_64_out_net_0[14]), .Y(
        SYN_3_0_a2_12_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \SYN_2_0_a2_13[0]  (.A(
        data_64_out_net_0[23]), .B(data_64_out_net_0[20]), .C(
        data_64_out_net_0[17]), .D(data_64_out_net_0[14]), .Y(
        SYN_2_0_a2_13_Z[0]));
    CFG4 #( .INIT(16'h6996) )  \SYN_0_a2_1_0[7]  (.A(
        data_64_out_net_0[12]), .B(data_64_out_net_0[59]), .C(
        data_64_out_net_0[35]), .D(data_64_out_net_0[61]), .Y(SYN_1[7])
        );
    CFG4 #( .INIT(16'h6996) )  \SYN_0_a2_12[7]  (.A(
        data_64_out_net_0[63]), .B(data_64_out_net_0[43]), .C(
        data_64_out_net_0[38]), .D(data_64_out_net_0[27]), .Y(
        SYN_0_a2_12_Z[7]));
    CFG4 #( .INIT(16'h6996) )  \SYN_0_a2_10[7]  (.A(SYN_6_3_Z[4]), .B(
        data_64_out_net_0[6]), .C(data_64_out_net_0[5]), .D(
        PF_TPSRAM_C0_0_R_DATA[7]), .Y(SYN_0_a2_10_Z[7]));
    CFG4 #( .INIT(16'h6996) )  \SYN_5_0_a2[3]  (.A(SYN_5_0_a2_16_Z[3]), 
        .B(SYN_5_0_a2_14_Z[3]), .C(SYN_5_0_a2_11_Z[3]), .D(
        SYN_5_0_a2_10_Z[3]), .Y(SYN_5[3]));
    CFG4 #( .INIT(16'h6996) )  \SYN_2_0_a2_9_0[0]  (.A(
        data_64_out_net_0[57]), .B(data_64_out_net_0[56]), .C(
        data_64_out_net_0[4]), .D(data_64_out_net_0[1]), .Y(
        SYN_2_0_a2_9[0]));
    CFG2 #( .INIT(4'h6) )  \SYN_4_0_a2_5[2]  (.A(data_64_out_net_0[20])
        , .B(data_64_out_net_0[21]), .Y(SYN_4_5[2]));
    CFG4 #( .INIT(16'h6996) )  \SYN_4_0_a2_15[2]  (.A(
        data_64_out_net_0[9]), .B(data_64_out_net_0[16]), .C(
        data_64_out_net_0[59]), .D(SYN_4_0_a2_10_Z[2]), .Y(
        SYN_4_0_a2_15_Z[2]));
    CFG4 #( .INIT(16'h6996) )  \SYN_8_0_a2_1_0[6]  (.A(
        data_64_out_net_0[61]), .B(data_64_out_net_0[53]), .C(
        data_64_out_net_0[35]), .D(data_64_out_net_0[27]), .Y(
        SYN_8_0_a2_1[6]));
    CFG3 #( .INIT(8'h96) )  \SYN_6_0[4]  (.A(data_64_out_net_0[49]), 
        .B(data_64_out_net_0[52]), .C(data_64_out_net_0[46]), .Y(
        SYN_6_0_Z[4]));
    CFG2 #( .INIT(4'h6) )  \SYN_3_0_a2_4[1]  (.A(data_64_out_net_0[25])
        , .B(data_64_out_net_0[32]), .Y(SYN_3_0_a2_4_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \SYN_7_0_a2_11[5]  (.A(
        SYN_7_0_a2_2_Z[5]), .B(data_64_out_net_0[53]), .C(
        data_64_out_net_0[27]), .D(N_27), .Y(SYN_7_0_a2_11_Z[5]));
    CFG2 #( .INIT(4'h6) )  \SYN_3_0_a2_5[1]  (.A(data_64_out_net_0[18])
        , .B(data_64_out_net_0[22]), .Y(SYN_3_5[1]));
    CFG4 #( .INIT(16'h6996) )  \SYN_6_13[4]  (.A(SYN_6_4_Z[4]), .B(
        SYN_6_3_0[4]), .C(data_64_out_net_0[36]), .D(
        data_64_out_net_0[35]), .Y(SYN_6_13_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \SYN_7_0_a2_12[5]  (.A(
        data_64_out_net_0[45]), .B(data_64_out_net_0[44]), .C(
        data_64_out_net_0[42]), .D(data_64_out_net_0[41]), .Y(
        SYN_7_0_a2_12_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \SYN_5_0_a2_7[3]  (.A(
        data_64_out_net_0[25]), .B(data_64_out_net_0[26]), .C(
        data_64_out_net_0[44]), .D(data_64_out_net_0[48]), .Y(
        SYN_5_0_a2_7_Z[3]));
    CFG4 #( .INIT(16'h6996) )  \SYN_0_a2_15[7]  (.A(SYN_0_a2_12_Z[7]), 
        .B(SYN_0_a2_3_Z[7]), .C(data_64_out_net_0[45]), .D(
        data_64_out_net_0[39]), .Y(SYN_0_a2_15_Z[7]));
    CFG4 #( .INIT(16'h6996) )  \SYN_0_a2[7]  (.A(SYN_0_a2_15_Z[7]), .B(
        SYN_0_a2_13_Z[7]), .C(SYN_0_a2_10_Z[7]), .D(SYN_0_a2_9_Z[7]), 
        .Y(SYN[7]));
    CFG2 #( .INIT(4'h6) )  \SYN_0_a2_8[7]  (.A(data_64_out_net_0[9]), 
        .B(data_64_out_net_0[16]), .Y(SYN_8[7]));
    CFG4 #( .INIT(16'h6996) )  \SYN_7_0_a2_6[5]  (.A(
        data_64_out_net_0[32]), .B(data_64_out_net_0[33]), .C(
        data_64_out_net_0[34]), .D(data_64_out_net_0[28]), .Y(
        SYN_7_0_a2_6_Z[5]));
    CFG3 #( .INIT(8'h96) )  \SYN_6_4[4]  (.A(data_64_out_net_0[34]), 
        .B(data_64_out_net_0[33]), .C(data_64_out_net_0[32]), .Y(
        SYN_6_4_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \SYN_4_0_a2_1[2]  (.A(
        data_64_out_net_0[3]), .B(data_64_out_net_0[29]), .C(
        data_64_out_net_0[19]), .D(data_64_out_net_0[40]), .Y(
        SYN_4_0_a2_1_Z[2]));
    CFG4 #( .INIT(16'h6996) )  \SYN_4_0_a2_12[2]  (.A(
        data_64_out_net_0[39]), .B(data_64_out_net_0[36]), .C(
        data_64_out_net_0[5]), .D(data_64_out_net_0[4]), .Y(
        SYN_4_0_a2_12_Z[2]));
    CFG4 #( .INIT(16'h6996) )  \SYN_3_0_a2_16[1]  (.A(
        SYN_3_0_a2_13_Z[1]), .B(SYN_3_0_a2_10_Z[1]), .C(
        SYN_3_0_a2_0_Z[1]), .D(data_64_out_net_0[60]), .Y(
        SYN_3_0_a2_16_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \SYN_2_0_a2_14[0]  (.A(
        data_64_out_net_0[47]), .B(data_64_out_net_0[24]), .C(
        data_64_out_net_0[7]), .D(data_64_out_net_0[6]), .Y(
        SYN_2_14[0]));
    CFG4 #( .INIT(16'h6996) )  \SYN_8_0_a2_10[6]  (.A(
        data_64_out_net_0[36]), .B(data_64_out_net_0[31]), .C(
        data_64_out_net_0[30]), .D(data_64_out_net_0[7]), .Y(
        SYN_8_0_a2_10_Z[6]));
    CFG4 #( .INIT(16'h6996) )  \SYN_3_0_a2_15[1]  (.A(
        SYN_3_0_a2_12_Z[1]), .B(SYN_3_0_a2_4_Z[1]), .C(
        data_64_out_net_0[31]), .D(data_64_out_net_0[1]), .Y(
        SYN_3_0_a2_15_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \SYN_3_0_a2_10[1]  (.A(
        data_64_out_net_0[54]), .B(data_64_out_net_0[51]), .C(
        data_64_out_net_0[11]), .D(data_64_out_net_0[8]), .Y(
        SYN_3_10[1]));
    CFG2 #( .INIT(4'h6) )  \SYN_6_12[4]  (.A(data_64_out_net_0[49]), 
        .B(data_64_out_net_0[52]), .Y(SYN_6_12_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \SYN_2_0_a2_12[0]  (.A(
        data_64_out_net_0[52]), .B(data_64_out_net_0[51]), .C(
        data_64_out_net_0[46]), .D(data_64_out_net_0[35]), .Y(
        SYN_2_0_a2_12_Z[0]));
    CFG2 #( .INIT(4'h6) )  \SYN_7_0_a2_0[5]  (.A(data_64_out_net_0[3]), 
        .B(data_64_out_net_0[29]), .Y(N_27));
    CFG4 #( .INIT(16'h6996) )  \SYN_4_0_a2_14[2]  (.A(
        data_64_out_net_0[63]), .B(data_64_out_net_0[62]), .C(
        data_64_out_net_0[43]), .D(data_64_out_net_0[26]), .Y(
        SYN_4_0_a2_14_Z[2]));
    CFG4 #( .INIT(16'h6996) )  \SYN_6_15[4]  (.A(SYN_6_0_Z[4]), .B(
        data_64_out_net_0[11]), .C(data_64_out_net_0[3]), .D(
        PF_TPSRAM_C0_0_R_DATA[4]), .Y(SYN_6_15_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \SYN_8_0_a2_9[6]  (.A(SYN_8_0_a2_1[6]), 
        .B(data_64_out_net_0[40]), .C(data_64_out_net_0[19]), .D(
        PF_TPSRAM_C0_0_R_DATA[6]), .Y(SYN_8_0_a2_9_Z[6]));
    CFG4 #( .INIT(16'h6996) )  \SYN_5_0_a2_16[3]  (.A(
        SYN_5_0_a2_12_Z[3]), .B(SYN_5_0_a2_7_Z[3]), .C(
        data_64_out_net_0[28]), .D(data_64_out_net_0[27]), .Y(
        SYN_5_0_a2_16_Z[3]));
    GND GND_Z (.Y(GND));
    VCC VCC_Z (.Y(VCC));
    CFG4 #( .INIT(16'h6996) )  \SYN_6_11[4]  (.A(data_64_out_net_0[45])
        , .B(data_64_out_net_0[42]), .C(data_64_out_net_0[39]), .D(
        data_64_out_net_0[37]), .Y(SYN_6_11_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \SYN_7_0_a2_2[5]  (.A(
        data_64_out_net_0[54]), .B(data_64_out_net_0[40]), .C(
        data_64_out_net_0[19]), .D(data_64_out_net_0[11]), .Y(
        SYN_7_0_a2_2_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \SYN_7_0_a2[5]  (.A(SYN_7_0_a2_16_Z[5]), 
        .B(SYN_7_0_a2_14_Z[5]), .C(SYN_7_0_a2_11_Z[5]), .D(
        SYN_7_0_a2_10_Z[5]), .Y(SYN_7[5]));
    CFG4 #( .INIT(16'h6996) )  \SYN_5_0_a2_10[3]  (.A(
        data_64_out_net_0[11]), .B(PF_TPSRAM_C0_0_R_DATA[3]), .C(N_31), 
        .D(N_27), .Y(SYN_5_0_a2_10_Z[3]));
    CFG4 #( .INIT(16'h6996) )  \SYN_4_0_a2_16[2]  (.A(
        SYN_4_0_a2_12_Z[2]), .B(SYN_4_0_a2_1_Z[2]), .C(
        data_64_out_net_0[17]), .D(data_64_out_net_0[10]), .Y(
        SYN_4_0_a2_16_Z[2]));
    CFG4 #( .INIT(16'hFFFE) )  ERRr (.A(SYN_2[0]), .B(SYN[7]), .C(
        ERRr_4_Z), .D(ERRr_2_Z), .Y(ERRr_c));
    CFG4 #( .INIT(16'h6996) )  \SYN_6_17[4]  (.A(SYN_6_13_Z[4]), .B(
        SYN_6_8_Z[4]), .C(SYN_4_5[2]), .D(data_64_out_net_0[24]), .Y(
        SYN_6_17_Z[4]));
    CFG4 #( .INIT(16'h6996) )  \SYN_7_0_a2_14[5]  (.A(
        data_64_out_net_0[63]), .B(data_64_out_net_0[60]), .C(
        data_64_out_net_0[47]), .D(data_64_out_net_0[46]), .Y(
        SYN_7_0_a2_14_Z[5]));
    CFG4 #( .INIT(16'h6996) )  \SYN_2_0_a2_0[0]  (.A(
        data_64_out_net_0[0]), .B(data_64_out_net_0[43]), .C(
        data_64_out_net_0[27]), .D(data_64_out_net_0[53]), .Y(
        SYN_2_0_a2_0_Z[0]));
    CFG3 #( .INIT(8'h96) )  \SYN_6_8[4]  (.A(data_64_out_net_0[15]), 
        .B(data_64_out_net_0[19]), .C(data_64_out_net_0[14]), .Y(
        SYN_6_8_Z[4]));
    CFG3 #( .INIT(8'h96) )  \SYN_3_0_a2_0[1]  (.A(data_64_out_net_0[0])
        , .B(data_64_out_net_0[43]), .C(SYN_1[7]), .Y(
        SYN_3_0_a2_0_Z[1]));
    CFG4 #( .INIT(16'h6996) )  \SYN_0_a2_13[7]  (.A(SYN_8[7]), .B(
        SYN_6[7]), .C(data_64_out_net_0[62]), .D(data_64_out_net_0[60])
        , .Y(SYN_0_a2_13_Z[7]));
    CFG2 #( .INIT(4'h6) )  \SYN_0_a2_6[7]  (.A(data_64_out_net_0[50]), 
        .B(data_64_out_net_0[58]), .Y(SYN_6[7]));
    CFG3 #( .INIT(8'h96) )  \SYN_0_a2_3[7]  (.A(data_64_out_net_0[57]), 
        .B(data_64_out_net_0[56]), .C(data_64_out_net_0[49]), .Y(
        SYN_0_a2_3_Z[7]));
    CFG4 #( .INIT(16'h6996) )  \SYN_5_0_a2_14[3]  (.A(SYN_2_14[0]), .B(
        data_64_out_net_0[51]), .C(data_64_out_net_0[41]), .D(
        data_64_out_net_0[38]), .Y(SYN_5_0_a2_14_Z[3]));
    CFG4 #( .INIT(16'h6996) )  \SYN_8_0_a2_13[6]  (.A(
        SYN_8_0_a2_9_Z[6]), .B(SYN_3_10[1]), .C(data_64_out_net_0[4]), 
        .D(data_64_out_net_0[1]), .Y(SYN_8_0_a2_13_Z[6]));
    CFG4 #( .INIT(16'h6996) )  \SYN_4_0_a2_13[2]  (.A(SYN_4_5[2]), .B(
        data_64_out_net_0[33]), .C(data_64_out_net_0[30]), .D(
        data_64_out_net_0[23]), .Y(SYN_4_0_a2_13_Z[2]));
    CFG4 #( .INIT(16'h6996) )  \SYN_8_0_a2_11[6]  (.A(SYN_6_12_Z[4]), 
        .B(data_64_out_net_0[62]), .C(data_64_out_net_0[55]), .D(
        data_64_out_net_0[42]), .Y(SYN_8_0_a2_11_Z[6]));
    CFG2 #( .INIT(4'h6) )  \SYN_7_0_a2_1[5]  (.A(data_64_out_net_0[0]), 
        .B(data_64_out_net_0[43]), .Y(N_32));
    CFG4 #( .INIT(16'h6996) )  \SYN_2_0_a2_11[0]  (.A(
        data_64_out_net_0[13]), .B(data_64_out_net_0[10]), .C(
        data_64_out_net_0[5]), .D(data_64_out_net_0[3]), .Y(
        SYN_2_0_a2_11_Z[0]));
    
endmodule


module de_v1(
       data_64_out_net_0,
       PF_TPSRAM_C0_0_R_DATA,
       ERRr_c
    );
input  [63:0] data_64_out_net_0;
input  [7:0] PF_TPSRAM_C0_0_R_DATA;
output ERRr_c;

    wire GND, VCC;
    
    de64_1 de1 (.PF_TPSRAM_C0_0_R_DATA({PF_TPSRAM_C0_0_R_DATA[7], 
        PF_TPSRAM_C0_0_R_DATA[6], PF_TPSRAM_C0_0_R_DATA[5], 
        PF_TPSRAM_C0_0_R_DATA[4], PF_TPSRAM_C0_0_R_DATA[3], 
        PF_TPSRAM_C0_0_R_DATA[2], PF_TPSRAM_C0_0_R_DATA[1], 
        PF_TPSRAM_C0_0_R_DATA[0]}), .data_64_out_net_0({
        data_64_out_net_0[63], data_64_out_net_0[62], 
        data_64_out_net_0[61], data_64_out_net_0[60], 
        data_64_out_net_0[59], data_64_out_net_0[58], 
        data_64_out_net_0[57], data_64_out_net_0[56], 
        data_64_out_net_0[55], data_64_out_net_0[54], 
        data_64_out_net_0[53], data_64_out_net_0[52], 
        data_64_out_net_0[51], data_64_out_net_0[50], 
        data_64_out_net_0[49], data_64_out_net_0[48], 
        data_64_out_net_0[47], data_64_out_net_0[46], 
        data_64_out_net_0[45], data_64_out_net_0[44], 
        data_64_out_net_0[43], data_64_out_net_0[42], 
        data_64_out_net_0[41], data_64_out_net_0[40], 
        data_64_out_net_0[39], data_64_out_net_0[38], 
        data_64_out_net_0[37], data_64_out_net_0[36], 
        data_64_out_net_0[35], data_64_out_net_0[34], 
        data_64_out_net_0[33], data_64_out_net_0[32], 
        data_64_out_net_0[31], data_64_out_net_0[30], 
        data_64_out_net_0[29], data_64_out_net_0[28], 
        data_64_out_net_0[27], data_64_out_net_0[26], 
        data_64_out_net_0[25], data_64_out_net_0[24], 
        data_64_out_net_0[23], data_64_out_net_0[22], 
        data_64_out_net_0[21], data_64_out_net_0[20], 
        data_64_out_net_0[19], data_64_out_net_0[18], 
        data_64_out_net_0[17], data_64_out_net_0[16], 
        data_64_out_net_0[15], data_64_out_net_0[14], 
        data_64_out_net_0[13], data_64_out_net_0[12], 
        data_64_out_net_0[11], data_64_out_net_0[10], 
        data_64_out_net_0[9], data_64_out_net_0[8], 
        data_64_out_net_0[7], data_64_out_net_0[6], 
        data_64_out_net_0[5], data_64_out_net_0[4], 
        data_64_out_net_0[3], data_64_out_net_0[2], 
        data_64_out_net_0[1], data_64_out_net_0[0]}), .ERRr_c(ERRr_c));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM(
       en64_RP2_0_OUTt,
       PF_TPSRAM_C0_0_R_DATA,
       W_ADDR_c,
       R_ADDR_c,
       W_EN_c,
       R_EN_c,
       CLK
    );
input  [7:0] en64_RP2_0_OUTt;
output [7:0] PF_TPSRAM_C0_0_R_DATA;
input  [13:0] W_ADDR_c;
input  [13:0] R_ADDR_c;
input  W_EN_c;
input  R_EN_c;
input  CLK;

    wire [19:1] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT;
    wire [19:0] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT;
    wire [19:1] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT;
    wire [19:0] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT;
    wire [19:1] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT;
    wire [19:0] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT;
    wire [19:1] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT;
    wire [19:0] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT;
    wire [19:1] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT;
    wire [19:0] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT;
    wire [19:1] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT;
    wire [19:0] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT;
    wire [19:1] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT;
    wire [19:0] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT;
    wire [19:1] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT;
    wire [19:0] PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT;
    wire VCC, GND, 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_SB_CORRECT, 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_DB_DETECT, 
        \Z\ACCESS_BUSY[0][4] , 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_SB_CORRECT, 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_DB_DETECT, 
        \Z\ACCESS_BUSY[0][3] , 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_SB_CORRECT, 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_DB_DETECT, 
        \Z\ACCESS_BUSY[0][6] , 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_SB_CORRECT, 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_DB_DETECT, 
        \Z\ACCESS_BUSY[0][0] , 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_SB_CORRECT, 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_DB_DETECT, 
        \Z\ACCESS_BUSY[0][7] , 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_SB_CORRECT, 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_DB_DETECT, 
        \Z\ACCESS_BUSY[0][1] , 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_SB_CORRECT, 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_DB_DETECT, 
        \Z\ACCESS_BUSY[0][5] , 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_SB_CORRECT, 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_DB_DETECT, 
        \Z\ACCESS_BUSY[0][2] ;
    
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_TPSRAM_C0_0%16384-16384%8-8%SPEED%0%4%TWO-PORT%ECC_EN-0")
         )  PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4 (.A_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_A_DOUT[1], 
        PF_TPSRAM_C0_0_R_DATA[4]}), .B_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[1], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_B_DOUT[0]}), 
        .DB_DETECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_DB_DETECT), 
        .SB_CORRECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C4_SB_CORRECT), 
        .ACCESS_BUSY(\Z\ACCESS_BUSY[0][4] ), .A_ADDR({R_ADDR_c[13], 
        R_ADDR_c[12], R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], 
        R_ADDR_c[8], R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], 
        R_ADDR_c[4], R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], 
        R_ADDR_c[0]}), .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .A_REN(R_EN_c), 
        .A_WEN({GND, GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[13], W_ADDR_c[12], 
        W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0]}), 
        .B_BLK_EN({W_EN_c, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, en64_RP2_0_OUTt[4]}), .B_REN(VCC), 
        .B_WEN({GND, VCC}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_TPSRAM_C0_0%16384-16384%8-8%SPEED%0%3%TWO-PORT%ECC_EN-0")
         )  PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3 (.A_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_A_DOUT[1], 
        PF_TPSRAM_C0_0_R_DATA[3]}), .B_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[1], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_B_DOUT[0]}), 
        .DB_DETECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_DB_DETECT), 
        .SB_CORRECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C3_SB_CORRECT), 
        .ACCESS_BUSY(\Z\ACCESS_BUSY[0][3] ), .A_ADDR({R_ADDR_c[13], 
        R_ADDR_c[12], R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], 
        R_ADDR_c[8], R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], 
        R_ADDR_c[4], R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], 
        R_ADDR_c[0]}), .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .A_REN(R_EN_c), 
        .A_WEN({GND, GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[13], W_ADDR_c[12], 
        W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0]}), 
        .B_BLK_EN({W_EN_c, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, en64_RP2_0_OUTt[3]}), .B_REN(VCC), 
        .B_WEN({GND, VCC}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    VCC VCC_Z (.Y(VCC));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_TPSRAM_C0_0%16384-16384%8-8%SPEED%0%1%TWO-PORT%ECC_EN-0")
         )  PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1 (.A_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_A_DOUT[1], 
        PF_TPSRAM_C0_0_R_DATA[1]}), .B_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[1], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_B_DOUT[0]}), 
        .DB_DETECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_DB_DETECT), 
        .SB_CORRECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C1_SB_CORRECT), 
        .ACCESS_BUSY(\Z\ACCESS_BUSY[0][1] ), .A_ADDR({R_ADDR_c[13], 
        R_ADDR_c[12], R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], 
        R_ADDR_c[8], R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], 
        R_ADDR_c[4], R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], 
        R_ADDR_c[0]}), .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .A_REN(R_EN_c), 
        .A_WEN({GND, GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[13], W_ADDR_c[12], 
        W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0]}), 
        .B_BLK_EN({W_EN_c, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, en64_RP2_0_OUTt[1]}), .B_REN(VCC), 
        .B_WEN({GND, VCC}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_TPSRAM_C0_0%16384-16384%8-8%SPEED%0%7%TWO-PORT%ECC_EN-0")
         )  PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7 (.A_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_A_DOUT[1], 
        PF_TPSRAM_C0_0_R_DATA[7]}), .B_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[1], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_B_DOUT[0]}), 
        .DB_DETECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_DB_DETECT), 
        .SB_CORRECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C7_SB_CORRECT), 
        .ACCESS_BUSY(\Z\ACCESS_BUSY[0][7] ), .A_ADDR({R_ADDR_c[13], 
        R_ADDR_c[12], R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], 
        R_ADDR_c[8], R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], 
        R_ADDR_c[4], R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], 
        R_ADDR_c[0]}), .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .A_REN(R_EN_c), 
        .A_WEN({GND, GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[13], W_ADDR_c[12], 
        W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0]}), 
        .B_BLK_EN({W_EN_c, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, en64_RP2_0_OUTt[7]}), .B_REN(VCC), 
        .B_WEN({GND, VCC}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_TPSRAM_C0_0%16384-16384%8-8%SPEED%0%6%TWO-PORT%ECC_EN-0")
         )  PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6 (.A_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_A_DOUT[1], 
        PF_TPSRAM_C0_0_R_DATA[6]}), .B_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[1], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_B_DOUT[0]}), 
        .DB_DETECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_DB_DETECT), 
        .SB_CORRECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C6_SB_CORRECT), 
        .ACCESS_BUSY(\Z\ACCESS_BUSY[0][6] ), .A_ADDR({R_ADDR_c[13], 
        R_ADDR_c[12], R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], 
        R_ADDR_c[8], R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], 
        R_ADDR_c[4], R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], 
        R_ADDR_c[0]}), .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .A_REN(R_EN_c), 
        .A_WEN({GND, GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[13], W_ADDR_c[12], 
        W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0]}), 
        .B_BLK_EN({W_EN_c, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, en64_RP2_0_OUTt[6]}), .B_REN(VCC), 
        .B_WEN({GND, VCC}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_TPSRAM_C0_0%16384-16384%8-8%SPEED%0%5%TWO-PORT%ECC_EN-0")
         )  PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5 (.A_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_A_DOUT[1], 
        PF_TPSRAM_C0_0_R_DATA[5]}), .B_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[1], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_B_DOUT[0]}), 
        .DB_DETECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_DB_DETECT), 
        .SB_CORRECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C5_SB_CORRECT), 
        .ACCESS_BUSY(\Z\ACCESS_BUSY[0][5] ), .A_ADDR({R_ADDR_c[13], 
        R_ADDR_c[12], R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], 
        R_ADDR_c[8], R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], 
        R_ADDR_c[4], R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], 
        R_ADDR_c[0]}), .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .A_REN(R_EN_c), 
        .A_WEN({GND, GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[13], W_ADDR_c[12], 
        W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0]}), 
        .B_BLK_EN({W_EN_c, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, en64_RP2_0_OUTt[5]}), .B_REN(VCC), 
        .B_WEN({GND, VCC}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_TPSRAM_C0_0%16384-16384%8-8%SPEED%0%2%TWO-PORT%ECC_EN-0")
         )  PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2 (.A_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_A_DOUT[1], 
        PF_TPSRAM_C0_0_R_DATA[2]}), .B_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[1], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_B_DOUT[0]}), 
        .DB_DETECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_DB_DETECT), 
        .SB_CORRECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C2_SB_CORRECT), 
        .ACCESS_BUSY(\Z\ACCESS_BUSY[0][2] ), .A_ADDR({R_ADDR_c[13], 
        R_ADDR_c[12], R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], 
        R_ADDR_c[8], R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], 
        R_ADDR_c[4], R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], 
        R_ADDR_c[0]}), .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .A_REN(R_EN_c), 
        .A_WEN({GND, GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[13], W_ADDR_c[12], 
        W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0]}), 
        .B_BLK_EN({W_EN_c, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, en64_RP2_0_OUTt[2]}), .B_REN(VCC), 
        .B_WEN({GND, VCC}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_TPSRAM_C0_0%16384-16384%8-8%SPEED%0%0%TWO-PORT%ECC_EN-0")
         )  PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0 (.A_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_A_DOUT[1], 
        PF_TPSRAM_C0_0_R_DATA[0]}), .B_DOUT({
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[19], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[18], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[17], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[16], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[15], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[14], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[13], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[12], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[11], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[10], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[9], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[8], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[7], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[6], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[5], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[4], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[3], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[2], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[1], 
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_B_DOUT[0]}), 
        .DB_DETECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_DB_DETECT), 
        .SB_CORRECT(
        PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM_R0C0_SB_CORRECT), 
        .ACCESS_BUSY(\Z\ACCESS_BUSY[0][0] ), .A_ADDR({R_ADDR_c[13], 
        R_ADDR_c[12], R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], 
        R_ADDR_c[8], R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], 
        R_ADDR_c[4], R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], 
        R_ADDR_c[0]}), .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .A_REN(R_EN_c), 
        .A_WEN({GND, GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[13], W_ADDR_c[12], 
        W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0]}), 
        .B_BLK_EN({W_EN_c, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, en64_RP2_0_OUTt[0]}), .B_REN(VCC), 
        .B_WEN({GND, VCC}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_TPSRAM_C0(
       R_ADDR_c,
       W_ADDR_c,
       PF_TPSRAM_C0_0_R_DATA,
       en64_RP2_0_OUTt,
       CLK,
       R_EN_c,
       W_EN_c
    );
input  [13:0] R_ADDR_c;
input  [13:0] W_ADDR_c;
output [7:0] PF_TPSRAM_C0_0_R_DATA;
input  [7:0] en64_RP2_0_OUTt;
input  CLK;
input  R_EN_c;
input  W_EN_c;

    wire GND, VCC;
    
    PF_TPSRAM_C0_PF_TPSRAM_C0_0_PF_TPSRAM PF_TPSRAM_C0_0 (
        .en64_RP2_0_OUTt({en64_RP2_0_OUTt[7], en64_RP2_0_OUTt[6], 
        en64_RP2_0_OUTt[5], en64_RP2_0_OUTt[4], en64_RP2_0_OUTt[3], 
        en64_RP2_0_OUTt[2], en64_RP2_0_OUTt[1], en64_RP2_0_OUTt[0]}), 
        .PF_TPSRAM_C0_0_R_DATA({PF_TPSRAM_C0_0_R_DATA[7], 
        PF_TPSRAM_C0_0_R_DATA[6], PF_TPSRAM_C0_0_R_DATA[5], 
        PF_TPSRAM_C0_0_R_DATA[4], PF_TPSRAM_C0_0_R_DATA[3], 
        PF_TPSRAM_C0_0_R_DATA[2], PF_TPSRAM_C0_0_R_DATA[1], 
        PF_TPSRAM_C0_0_R_DATA[0]}), .W_ADDR_c({W_ADDR_c[13], 
        W_ADDR_c[12], W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], 
        W_ADDR_c[8], W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], 
        W_ADDR_c[4], W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], 
        W_ADDR_c[0]}), .R_ADDR_c({R_ADDR_c[13], R_ADDR_c[12], 
        R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0]}), .W_EN_c(
        W_EN_c), .R_EN_c(R_EN_c), .CLK(CLK));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module error_gen(
       data_64_out_net_0,
       R_DATA_c,
       selectt_c
    );
output [63:0] data_64_out_net_0;
input  [77:0] R_DATA_c;
input  [63:0] selectt_c;

    wire [63:63] OUTt_0_iv_0_o2_5_42_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_41_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_40_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_39_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_38_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_37_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_36_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_35_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_34_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_33_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_32_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_31_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_30_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_29_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_53_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_52_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_51_Z;
    wire [63:63] OUTt_0_iv_0_o2_5_50_Z;
    wire N_206, N_205, N_204, N_203, N_202, N_201, N_200, N_199, N_196, 
        N_210, N_209, N_208, N_207, GND, VCC;
    
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI21ED1[54]  (.A(N_210), .B(N_203)
        , .C(N_199), .D(R_DATA_c[66]), .Y(data_64_out_net_0[54]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIOG7D1[22]  (.A(N_208), .B(N_203)
        , .C(N_199), .D(R_DATA_c[26]), .Y(data_64_out_net_0[22]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI79K11[46]  (.A(N_210), .B(N_205)
        , .C(N_200), .D(R_DATA_c[56]), .Y(data_64_out_net_0[46]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIMFC91[17]  (.A(N_207), .B(N_204)
        , .C(N_202), .D(R_DATA_c[21]), .Y(data_64_out_net_0[17]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI188V[5]  (.A(N_207), .B(N_205), 
        .C(N_204), .D(R_DATA_c[5]), .Y(data_64_out_net_0[5]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_34[63]  (.A(
        selectt_c[45]), .B(selectt_c[44]), .C(selectt_c[43]), .D(
        selectt_c[42]), .Y(OUTt_0_iv_0_o2_5_34_Z[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNINID11[11]  (.A(N_207), .B(N_206)
        , .C(N_200), .D(R_DATA_c[13]), .Y(data_64_out_net_0[11]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI2PV41[51]  (.A(N_209), .B(N_203)
        , .C(N_202), .D(R_DATA_c[63]), .Y(data_64_out_net_0[51]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_41[63]  (.A(
        selectt_c[25]), .B(selectt_c[24]), .C(selectt_c[23]), .D(
        selectt_c[22]), .Y(OUTt_0_iv_0_o2_5_41_Z[63]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_40[63]  (.A(
        selectt_c[21]), .B(selectt_c[20]), .C(selectt_c[19]), .D(
        selectt_c[18]), .Y(OUTt_0_iv_0_o2_5_40_Z[63]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_33[63]  (.A(
        selectt_c[41]), .B(selectt_c[40]), .C(selectt_c[39]), .D(
        selectt_c[38]), .Y(OUTt_0_iv_0_o2_5_33_Z[63]));
    CFG2 #( .INIT(4'h7) )  \OUTt_0_iv_0_o2_3[63]  (.A(selectt_c[2]), 
        .B(selectt_c[4]), .Y(N_199));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIT38V[3]  (.A(N_207), .B(N_206), 
        .C(N_203), .D(R_DATA_c[3]), .Y(data_64_out_net_0[3]));
    CFG2 #( .INIT(4'hB) )  \OUTt_0_iv_i_o2_1[41]  (.A(selectt_c[1]), 
        .B(selectt_c[3]), .Y(N_201));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIOEV41[41]  (.A(N_209), .B(N_206)
        , .C(N_201), .D(R_DATA_c[51]), .Y(data_64_out_net_0[41]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_31[63]  (.A(
        selectt_c[33]), .B(selectt_c[32]), .C(selectt_c[15]), .D(
        selectt_c[14]), .Y(OUTt_0_iv_0_o2_5_31_Z[63]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_30[63]  (.A(
        selectt_c[13]), .B(selectt_c[12]), .C(selectt_c[11]), .D(
        selectt_c[10]), .Y(OUTt_0_iv_0_o2_5_30_Z[63]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_38[63]  (.A(
        selectt_c[61]), .B(selectt_c[60]), .C(selectt_c[59]), .D(
        selectt_c[58]), .Y(OUTt_0_iv_0_o2_5_38_Z[63]));
    CFG2 #( .INIT(4'hE) )  \OUTt_0_iv_i_o2_1[43]  (.A(selectt_c[2]), 
        .B(selectt_c[4]), .Y(N_206));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI089V[9]  (.A(N_207), .B(N_206), 
        .C(N_201), .D(R_DATA_c[11]), .Y(data_64_out_net_0[9]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNITRH91[38]  (.A(N_210), .B(N_205)
        , .C(N_203), .D(R_DATA_c[46]), .Y(data_64_out_net_0[38]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIKC7D1[20]  (.A(N_208), .B(N_204)
        , .C(N_199), .D(R_DATA_c[24]), .Y(data_64_out_net_0[20]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIUIT41[35]  (.A(N_209), .B(N_206)
        , .C(N_203), .D(R_DATA_c[43]), .Y(data_64_out_net_0[35]));
    CFG3 #( .INIT(8'hF7) )  \OUTt_0_iv_0_o2_0[63]  (.A(selectt_c[5]), 
        .B(selectt_c[0]), .C(N_196), .Y(N_209));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI0NV41[45]  (.A(N_209), .B(N_205)
        , .C(N_201), .D(R_DATA_c[55]), .Y(data_64_out_net_0[45]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI7TU41[49]  (.A(N_209), .B(N_204)
        , .C(N_202), .D(R_DATA_c[61]), .Y(data_64_out_net_0[49]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_29[63]  (.A(
        selectt_c[9]), .B(selectt_c[8]), .C(selectt_c[7]), .D(
        selectt_c[6]), .Y(OUTt_0_iv_0_o2_5_29_Z[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIOHC91[18]  (.A(N_208), .B(N_203)
        , .C(N_202), .D(R_DATA_c[22]), .Y(data_64_out_net_0[18]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI5SR81[61]  (.A(N_209), .B(N_201)
        , .C(N_199), .D(R_DATA_c[75]), .Y(data_64_out_net_0[61]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNICFL11[58]  (.A(N_210), .B(N_202)
        , .C(N_200), .D(R_DATA_c[72]), .Y(data_64_out_net_0[58]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIPNH91[36]  (.A(N_210), .B(N_205)
        , .C(N_204), .D(R_DATA_c[44]), .Y(data_64_out_net_0[36]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIV58V[4]  (.A(N_208), .B(N_205), 
        .C(N_204), .D(R_DATA_c[4]), .Y(data_64_out_net_0[4]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNITM8D1[29]  (.A(N_207), .B(N_201)
        , .C(N_199), .D(R_DATA_c[35]), .Y(data_64_out_net_0[29]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNILJH91[34]  (.A(N_210), .B(N_206)
        , .C(N_203), .D(R_DATA_c[42]), .Y(data_64_out_net_0[34]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIKFE91[25]  (.A(N_207), .B(N_202)
        , .C(N_201), .D(R_DATA_c[31]), .Y(data_64_out_net_0[25]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_37[63]  (.A(
        selectt_c[57]), .B(selectt_c[56]), .C(selectt_c[55]), .D(
        selectt_c[54]), .Y(OUTt_0_iv_0_o2_5_37_Z[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNILDS01[63]  (.A(N_209), .B(N_200)
        , .C(N_199), .D(R_DATA_c[77]), .Y(data_64_out_net_0[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNICEG51[62]  (.A(N_210), .B(N_200)
        , .C(N_199), .D(R_DATA_c[76]), .Y(data_64_out_net_0[62]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_35[63]  (.A(
        selectt_c[49]), .B(selectt_c[48]), .C(selectt_c[47]), .D(
        selectt_c[46]), .Y(OUTt_0_iv_0_o2_5_35_Z[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIKDC91[16]  (.A(N_208), .B(N_204)
        , .C(N_202), .D(R_DATA_c[20]), .Y(data_64_out_net_0[16]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIIDE91[24]  (.A(N_208), .B(N_202)
        , .C(N_201), .D(R_DATA_c[30]), .Y(data_64_out_net_0[24]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNISTK91[56]  (.A(N_210), .B(N_202)
        , .C(N_201), .D(R_DATA_c[70]), .Y(data_64_out_net_0[56]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIG80T[47]  (.A(N_209), .B(N_205), 
        .C(N_200), .D(R_DATA_c[57]), .Y(data_64_out_net_0[47]));
    CFG2 #( .INIT(4'hD) )  \OUTt_0_iv_i_o2_1[35]  (.A(selectt_c[1]), 
        .B(selectt_c[3]), .Y(N_203));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIPV7V[1]  (.A(N_207), .B(N_206), 
        .C(N_204), .D(R_DATA_c[1]), .Y(data_64_out_net_0[1]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI5C8V[7]  (.A(N_207), .B(N_205), 
        .C(N_203), .D(R_DATA_c[7]), .Y(data_64_out_net_0[7]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIRK8D1[28]  (.A(N_208), .B(N_201)
        , .C(N_199), .D(R_DATA_c[34]), .Y(data_64_out_net_0[28]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_39[63]  (.A(
        selectt_c[63]), .B(selectt_c[62]), .C(selectt_c[17]), .D(
        selectt_c[16]), .Y(OUTt_0_iv_0_o2_5_39_Z[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIUSDD1[52]  (.A(N_210), .B(N_204)
        , .C(N_199), .D(R_DATA_c[64]), .Y(data_64_out_net_0[52]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI41F11[27]  (.A(N_207), .B(N_202)
        , .C(N_200), .D(R_DATA_c[33]), .Y(data_64_out_net_0[27]));
    CFG3 #( .INIT(8'hFB) )  \OUTt_0_iv_i_o2_0[31]  (.A(selectt_c[5]), 
        .B(selectt_c[0]), .C(N_196), .Y(N_207));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI3A8V[6]  (.A(N_208), .B(N_205), 
        .C(N_203), .D(R_DATA_c[6]), .Y(data_64_out_net_0[6]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNISSFD1[60]  (.A(N_210), .B(N_201)
        , .C(N_199), .D(R_DATA_c[74]), .Y(data_64_out_net_0[60]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNID7D91[12]  (.A(N_208), .B(N_205)
        , .C(N_201), .D(R_DATA_c[14]), .Y(data_64_out_net_0[12]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_36[63]  (.A(
        selectt_c[53]), .B(selectt_c[52]), .C(selectt_c[51]), .D(
        selectt_c[50]), .Y(OUTt_0_iv_0_o2_5_36_Z[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIU59V[8]  (.A(N_208), .B(N_206), 
        .C(N_201), .D(R_DATA_c[10]), .Y(data_64_out_net_0[8]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI5T051[57]  (.A(N_209), .B(N_202)
        , .C(N_201), .D(R_DATA_c[71]), .Y(data_64_out_net_0[57]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI7SP81[53]  (.A(N_209), .B(N_204)
        , .C(N_199), .D(R_DATA_c[65]), .Y(data_64_out_net_0[53]));
    CFG2 #( .INIT(4'hB) )  \OUTt_0_iv_i_o2_1[49]  (.A(selectt_c[2]), 
        .B(selectt_c[4]), .Y(N_202));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIVQD11[15]  (.A(N_207), .B(N_205)
        , .C(N_200), .D(R_DATA_c[17]), .Y(data_64_out_net_0[15]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIPPJ91[50]  (.A(N_210), .B(N_203)
        , .C(N_202), .D(R_DATA_c[62]), .Y(data_64_out_net_0[50]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI6RT41[39]  (.A(N_209), .B(N_205)
        , .C(N_203), .D(R_DATA_c[47]), .Y(data_64_out_net_0[39]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIQET41[33]  (.A(N_209), .B(N_206)
        , .C(N_204), .D(R_DATA_c[41]), .Y(data_64_out_net_0[33]));
    GND GND_Z (.Y(GND));
    VCC VCC_Z (.Y(VCC));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIME7D1[21]  (.A(N_207), .B(N_204)
        , .C(N_199), .D(R_DATA_c[25]), .Y(data_64_out_net_0[21]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNINNJ91[44]  (.A(N_210), .B(N_205)
        , .C(N_201), .D(R_DATA_c[54]), .Y(data_64_out_net_0[44]));
    CFG3 #( .INIT(8'hFE) )  \OUTt_0_iv_i_o2_0[30]  (.A(selectt_c[5]), 
        .B(selectt_c[0]), .C(N_196), .Y(N_208));
    CFG2 #( .INIT(4'h7) )  \OUTt_0_iv_0_o2_4[63]  (.A(selectt_c[1]), 
        .B(selectt_c[3]), .Y(N_200));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNILE1T[59]  (.A(N_209), .B(N_202), 
        .C(N_200), .D(R_DATA_c[73]), .Y(data_64_out_net_0[59]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIFFJ91[40]  (.A(N_210), .B(N_206)
        , .C(N_201), .D(R_DATA_c[50]), .Y(data_64_out_net_0[40]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIB0Q81[55]  (.A(N_209), .B(N_203)
        , .C(N_199), .D(R_DATA_c[67]), .Y(data_64_out_net_0[55]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI2U951[30]  (.A(N_208), .B(N_200)
        , .C(N_199), .D(R_DATA_c[36]), .Y(data_64_out_net_0[30]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNILGD11[10]  (.A(N_208), .B(N_206)
        , .C(N_200), .D(R_DATA_c[12]), .Y(data_64_out_net_0[10]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_52[63]  (.A(
        OUTt_0_iv_0_o2_5_37_Z[63]), .B(OUTt_0_iv_0_o2_5_36_Z[63]), .C(
        OUTt_0_iv_0_o2_5_35_Z[63]), .D(OUTt_0_iv_0_o2_5_34_Z[63]), .Y(
        OUTt_0_iv_0_o2_5_52_Z[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNITOD11[14]  (.A(N_208), .B(N_205)
        , .C(N_200), .D(R_DATA_c[16]), .Y(data_64_out_net_0[14]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI800T[43]  (.A(N_209), .B(N_206), 
        .C(N_200), .D(R_DATA_c[53]), .Y(data_64_out_net_0[43]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5[63]  (.A(
        OUTt_0_iv_0_o2_5_53_Z[63]), .B(OUTt_0_iv_0_o2_5_52_Z[63]), .C(
        OUTt_0_iv_0_o2_5_51_Z[63]), .D(OUTt_0_iv_0_o2_5_50_Z[63]), .Y(
        N_196));
    CFG2 #( .INIT(4'hD) )  \OUTt_0_iv_i_o2_1[47]  (.A(selectt_c[2]), 
        .B(selectt_c[4]), .Y(N_205));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIF9D91[13]  (.A(N_207), .B(N_205)
        , .C(N_201), .D(R_DATA_c[15]), .Y(data_64_out_net_0[13]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI2VE11[26]  (.A(N_208), .B(N_202)
        , .C(N_200), .D(R_DATA_c[32]), .Y(data_64_out_net_0[26]));
    CFG3 #( .INIT(8'hFD) )  \OUTt_0_iv_i_o2_0[62]  (.A(selectt_c[5]), 
        .B(selectt_c[0]), .C(N_196), .Y(N_210));
    CFG2 #( .INIT(4'hE) )  \OUTt_0_iv_i_o2_1[33]  (.A(selectt_c[1]), 
        .B(selectt_c[3]), .Y(N_204));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_53[63]  (.A(
        OUTt_0_iv_0_o2_5_41_Z[63]), .B(OUTt_0_iv_0_o2_5_40_Z[63]), .C(
        OUTt_0_iv_0_o2_5_39_Z[63]), .D(OUTt_0_iv_0_o2_5_38_Z[63]), .Y(
        OUTt_0_iv_0_o2_5_53_Z[63]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_42[63]  (.A(
        selectt_c[29]), .B(selectt_c[28]), .C(selectt_c[27]), .D(
        selectt_c[26]), .Y(OUTt_0_iv_0_o2_5_42_Z[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIQJC91[19]  (.A(N_207), .B(N_203)
        , .C(N_202), .D(R_DATA_c[23]), .Y(data_64_out_net_0[19]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIUTI91[48]  (.A(N_210), .B(N_204)
        , .C(N_202), .D(R_DATA_c[60]), .Y(data_64_out_net_0[48]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI40A51[31]  (.A(N_207), .B(N_200)
        , .C(N_199), .D(R_DATA_c[37]), .Y(data_64_out_net_0[31]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_51[63]  (.A(
        OUTt_0_iv_0_o2_5_33_Z[63]), .B(OUTt_0_iv_0_o2_5_32_Z[63]), .C(
        OUTt_0_iv_0_o2_5_31_Z[63]), .D(OUTt_0_iv_0_o2_5_30_Z[63]), .Y(
        OUTt_0_iv_0_o2_5_51_Z[63]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_50[63]  (.A(
        selectt_c[31]), .B(selectt_c[30]), .C(
        OUTt_0_iv_0_o2_5_42_Z[63]), .D(OUTt_0_iv_0_o2_5_29_Z[63]), .Y(
        OUTt_0_iv_0_o2_5_50_Z[63]));
    CFG4 #( .INIT(16'hFFFE) )  \OUTt_0_iv_0_o2_5_32[63]  (.A(
        selectt_c[37]), .B(selectt_c[36]), .C(selectt_c[35]), .D(
        selectt_c[34]), .Y(OUTt_0_iv_0_o2_5_32_Z[63]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIHFH91[32]  (.A(N_210), .B(N_206)
        , .C(N_204), .D(R_DATA_c[40]), .Y(data_64_out_net_0[32]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNI2NT41[37]  (.A(N_209), .B(N_205)
        , .C(N_204), .D(R_DATA_c[45]), .Y(data_64_out_net_0[37]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIV0K11[42]  (.A(N_210), .B(N_206)
        , .C(N_200), .D(R_DATA_c[52]), .Y(data_64_out_net_0[42]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIR18V[2]  (.A(N_208), .B(N_206), 
        .C(N_203), .D(R_DATA_c[2]), .Y(data_64_out_net_0[2]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNIQI7D1[23]  (.A(N_207), .B(N_203)
        , .C(N_199), .D(R_DATA_c[27]), .Y(data_64_out_net_0[23]));
    CFG4 #( .INIT(16'hFE01) )  \INn_RNINT7V[0]  (.A(N_208), .B(N_206), 
        .C(N_204), .D(R_DATA_c[0]), .Y(data_64_out_net_0[0]));
    
endmodule


module PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM(
       R_DATA_c,
       WBYTE_EN_c,
       W_DATA_c,
       W_ADDR_c,
       R_ADDR_c,
       CLK,
       R_EN_c,
       W_EN_c
    );
output [79:0] R_DATA_c;
input  [7:0] WBYTE_EN_c;
input  [79:0] W_DATA_c;
input  [13:0] W_ADDR_c;
input  [13:0] R_ADDR_c;
input  CLK;
input  R_EN_c;
input  W_EN_c;

    wire CFG2_7_Y, \Z\BLKX2[2] , CFG2_4_Y, CFG2_3_Y, \Z\BLKY2[4] , 
        CFG2_6_Y, \Z\BLKY2[1] , CFG2_0_Y, CFG2_5_Y, \Z\BLKY2[3] , 
        \Z\BLKX2[0] , \Z\BLKY2[5] , \Z\BLKY2[7] , CFG2_1_Y, 
        \Z\BLKY2[6] , CFG2_2_Y, \Z\BLKY2[2] , \Z\BLKX2[4] , 
        \Z\BLKX2[1] , \Z\BLKX2[3] , \Z\BLKX2[5] , \Z\BLKX2[7] , 
        \Z\BLKY2[0] , \Z\BLKX2[6] , OR4_303_Y, \Z\R_DATA_TEMPR28[28] , 
        \Z\R_DATA_TEMPR29[28] , \Z\R_DATA_TEMPR30[28] , 
        \Z\R_DATA_TEMPR31[28] , OR4_169_Y, \Z\R_DATA_TEMPR8[78] , 
        \Z\R_DATA_TEMPR9[78] , \Z\R_DATA_TEMPR10[78] , 
        \Z\R_DATA_TEMPR11[78] , OR2_25_Y, \Z\R_DATA_TEMPR20[30] , 
        \Z\R_DATA_TEMPR21[30] , OR4_130_Y, \Z\R_DATA_TEMPR16[35] , 
        \Z\R_DATA_TEMPR17[35] , \Z\R_DATA_TEMPR18[35] , 
        \Z\R_DATA_TEMPR19[35] , OR4_337_Y, \Z\R_DATA_TEMPR8[71] , 
        \Z\R_DATA_TEMPR9[71] , \Z\R_DATA_TEMPR10[71] , 
        \Z\R_DATA_TEMPR11[71] , OR4_615_Y, \Z\R_DATA_TEMPR8[75] , 
        \Z\R_DATA_TEMPR9[75] , \Z\R_DATA_TEMPR10[75] , 
        \Z\R_DATA_TEMPR11[75] , OR4_321_Y, \Z\R_DATA_TEMPR0[5] , 
        \Z\R_DATA_TEMPR1[5] , \Z\R_DATA_TEMPR2[5] , 
        \Z\R_DATA_TEMPR3[5] , OR4_98_Y, \Z\R_DATA_TEMPR8[27] , 
        \Z\R_DATA_TEMPR9[27] , \Z\R_DATA_TEMPR10[27] , 
        \Z\R_DATA_TEMPR11[27] , OR4_630_Y, OR4_511_Y, OR4_666_Y, 
        OR4_20_Y, OR4_550_Y, OR4_712_Y, OR4_238_Y, OR4_75_Y, OR4_64_Y, 
        OR4_514_Y, OR4_368_Y, \Z\R_DATA_TEMPR4[11] , 
        \Z\R_DATA_TEMPR5[11] , \Z\R_DATA_TEMPR6[11] , 
        \Z\R_DATA_TEMPR7[11] , OR4_633_Y, OR4_536_Y, OR4_217_Y, 
        OR4_524_Y, \Z\R_DATA_TEMPR0[19] , \Z\R_DATA_TEMPR1[19] , 
        \Z\R_DATA_TEMPR2[19] , \Z\R_DATA_TEMPR3[19] , OR4_570_Y, 
        \Z\R_DATA_TEMPR16[42] , \Z\R_DATA_TEMPR17[42] , 
        \Z\R_DATA_TEMPR18[42] , \Z\R_DATA_TEMPR19[42] , OR4_579_Y, 
        \Z\R_DATA_TEMPR12[26] , \Z\R_DATA_TEMPR13[26] , 
        \Z\R_DATA_TEMPR14[26] , \Z\R_DATA_TEMPR15[26] , OR4_47_Y, 
        \Z\R_DATA_TEMPR12[34] , \Z\R_DATA_TEMPR13[34] , 
        \Z\R_DATA_TEMPR14[34] , \Z\R_DATA_TEMPR15[34] , OR4_500_Y, 
        \Z\R_DATA_TEMPR12[58] , \Z\R_DATA_TEMPR13[58] , 
        \Z\R_DATA_TEMPR14[58] , \Z\R_DATA_TEMPR15[58] , OR4_166_Y, 
        \Z\R_DATA_TEMPR4[34] , \Z\R_DATA_TEMPR5[34] , 
        \Z\R_DATA_TEMPR6[34] , \Z\R_DATA_TEMPR7[34] , OR4_509_Y, 
        \Z\R_DATA_TEMPR8[16] , \Z\R_DATA_TEMPR9[16] , 
        \Z\R_DATA_TEMPR10[16] , \Z\R_DATA_TEMPR11[16] , GND, 
        \Z\BLKY1[0] , \Z\R_DATA_TEMPR5[20] , \Z\R_DATA_TEMPR5[21] , 
        \Z\R_DATA_TEMPR5[22] , \Z\R_DATA_TEMPR5[23] , 
        \Z\R_DATA_TEMPR5[24] , \Z\R_DATA_TEMPR5[25] , 
        \Z\R_DATA_TEMPR5[26] , \Z\R_DATA_TEMPR5[27] , 
        \Z\R_DATA_TEMPR5[28] , \Z\R_DATA_TEMPR5[29] , 
        \Z\R_DATA_TEMPR5[30] , \Z\R_DATA_TEMPR5[31] , 
        \Z\R_DATA_TEMPR5[32] , \Z\R_DATA_TEMPR5[33] , 
        \Z\R_DATA_TEMPR5[35] , \Z\R_DATA_TEMPR5[36] , 
        \Z\R_DATA_TEMPR5[37] , \Z\R_DATA_TEMPR5[38] , 
        \Z\R_DATA_TEMPR5[39] , VCC, \Z\BLKX1[0] , \Z\R_DATA_TEMPR5[0] , 
        \Z\R_DATA_TEMPR5[1] , \Z\R_DATA_TEMPR5[2] , 
        \Z\R_DATA_TEMPR5[3] , \Z\R_DATA_TEMPR5[4] , 
        \Z\R_DATA_TEMPR5[5] , \Z\R_DATA_TEMPR5[6] , 
        \Z\R_DATA_TEMPR5[7] , \Z\R_DATA_TEMPR5[8] , 
        \Z\R_DATA_TEMPR5[9] , \Z\R_DATA_TEMPR5[10] , 
        \Z\R_DATA_TEMPR5[12] , \Z\R_DATA_TEMPR5[13] , 
        \Z\R_DATA_TEMPR5[14] , \Z\R_DATA_TEMPR5[15] , 
        \Z\R_DATA_TEMPR5[16] , \Z\R_DATA_TEMPR5[17] , 
        \Z\R_DATA_TEMPR5[18] , \Z\R_DATA_TEMPR5[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0_DB_DETECT, 
        \Z\ACCESS_BUSY[5][0] , OR4_40_Y, \Z\R_DATA_TEMPR4[19] , 
        \Z\R_DATA_TEMPR6[19] , \Z\R_DATA_TEMPR7[19] , OR4_490_Y, 
        \Z\R_DATA_TEMPR16[2] , \Z\R_DATA_TEMPR17[2] , 
        \Z\R_DATA_TEMPR18[2] , \Z\R_DATA_TEMPR19[2] , OR4_315_Y, 
        \Z\R_DATA_TEMPR28[24] , \Z\R_DATA_TEMPR29[24] , 
        \Z\R_DATA_TEMPR30[24] , \Z\R_DATA_TEMPR31[24] , OR2_5_Y, 
        \Z\R_DATA_TEMPR20[40] , \Z\R_DATA_TEMPR21[40] , OR4_469_Y, 
        OR4_333_Y, OR2_34_Y, \Z\R_DATA_TEMPR22[63] , 
        \Z\R_DATA_TEMPR23[63] , OR4_686_Y, OR4_572_Y, OR4_718_Y, 
        OR4_71_Y, OR4_610_Y, OR4_522_Y, \Z\R_DATA_TEMPR12[42] , 
        \Z\R_DATA_TEMPR13[42] , \Z\R_DATA_TEMPR14[42] , 
        \Z\R_DATA_TEMPR15[42] , OR4_635_Y, OR4_110_Y, OR2_56_Y, 
        \Z\R_DATA_TEMPR22[21] , \Z\R_DATA_TEMPR23[21] , OR4_462_Y, 
        OR4_596_Y, OR4_297_Y, OR4_445_Y, OR4_80_Y, OR4_61_Y, 
        \Z\R_DATA_TEMPR0[59] , \Z\R_DATA_TEMPR1[59] , 
        \Z\R_DATA_TEMPR2[59] , \Z\R_DATA_TEMPR3[59] , OR4_644_Y, 
        \Z\R_DATA_TEMPR4[36] , \Z\R_DATA_TEMPR6[36] , 
        \Z\R_DATA_TEMPR7[36] , OR4_391_Y, \Z\R_DATA_TEMPR24[33] , 
        \Z\R_DATA_TEMPR25[33] , \Z\R_DATA_TEMPR26[33] , 
        \Z\R_DATA_TEMPR27[33] , OR4_478_Y, \Z\R_DATA_TEMPR8[2] , 
        \Z\R_DATA_TEMPR9[2] , \Z\R_DATA_TEMPR10[2] , 
        \Z\R_DATA_TEMPR11[2] , OR4_363_Y, \Z\R_DATA_TEMPR12[62] , 
        \Z\R_DATA_TEMPR13[62] , \Z\R_DATA_TEMPR14[62] , 
        \Z\R_DATA_TEMPR15[62] , OR4_471_Y, \Z\R_DATA_TEMPR4[16] , 
        \Z\R_DATA_TEMPR6[16] , \Z\R_DATA_TEMPR7[16] , OR4_408_Y, 
        \Z\R_DATA_TEMPR16[62] , \Z\R_DATA_TEMPR17[62] , 
        \Z\R_DATA_TEMPR18[62] , \Z\R_DATA_TEMPR19[62] , OR4_74_Y, 
        \Z\R_DATA_TEMPR16[20] , \Z\R_DATA_TEMPR17[20] , 
        \Z\R_DATA_TEMPR18[20] , \Z\R_DATA_TEMPR19[20] , OR4_249_Y, 
        OR4_133_Y, OR4_532_Y, OR4_634_Y, OR4_401_Y, 
        \Z\R_DATA_TEMPR24[56] , \Z\R_DATA_TEMPR25[56] , 
        \Z\R_DATA_TEMPR26[56] , \Z\R_DATA_TEMPR27[56] , OR4_221_Y, 
        \Z\R_DATA_TEMPR4[39] , \Z\R_DATA_TEMPR6[39] , 
        \Z\R_DATA_TEMPR7[39] , OR4_246_Y, \Z\R_DATA_TEMPR24[4] , 
        \Z\R_DATA_TEMPR25[4] , \Z\R_DATA_TEMPR26[4] , 
        \Z\R_DATA_TEMPR27[4] , \Z\BLKY0[0] , \Z\R_DATA_TEMPR10[20] , 
        \Z\R_DATA_TEMPR10[21] , \Z\R_DATA_TEMPR10[22] , 
        \Z\R_DATA_TEMPR10[23] , \Z\R_DATA_TEMPR10[24] , 
        \Z\R_DATA_TEMPR10[25] , \Z\R_DATA_TEMPR10[26] , 
        \Z\R_DATA_TEMPR10[28] , \Z\R_DATA_TEMPR10[29] , 
        \Z\R_DATA_TEMPR10[30] , \Z\R_DATA_TEMPR10[31] , 
        \Z\R_DATA_TEMPR10[32] , \Z\R_DATA_TEMPR10[33] , 
        \Z\R_DATA_TEMPR10[34] , \Z\R_DATA_TEMPR10[35] , 
        \Z\R_DATA_TEMPR10[36] , \Z\R_DATA_TEMPR10[37] , 
        \Z\R_DATA_TEMPR10[38] , \Z\R_DATA_TEMPR10[39] , \Z\BLKX0[0] , 
        \Z\R_DATA_TEMPR10[0] , \Z\R_DATA_TEMPR10[1] , 
        \Z\R_DATA_TEMPR10[3] , \Z\R_DATA_TEMPR10[4] , 
        \Z\R_DATA_TEMPR10[5] , \Z\R_DATA_TEMPR10[6] , 
        \Z\R_DATA_TEMPR10[7] , \Z\R_DATA_TEMPR10[8] , 
        \Z\R_DATA_TEMPR10[9] , \Z\R_DATA_TEMPR10[10] , 
        \Z\R_DATA_TEMPR10[11] , \Z\R_DATA_TEMPR10[12] , 
        \Z\R_DATA_TEMPR10[13] , \Z\R_DATA_TEMPR10[14] , 
        \Z\R_DATA_TEMPR10[15] , \Z\R_DATA_TEMPR10[17] , 
        \Z\R_DATA_TEMPR10[18] , \Z\R_DATA_TEMPR10[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0_DB_DETECT, 
        \Z\ACCESS_BUSY[10][0] , OR4_214_Y, OR4_306_Y, 
        \Z\R_DATA_TEMPR22[30] , \Z\R_DATA_TEMPR23[30] , OR4_553_Y, 
        \Z\R_DATA_TEMPR16[46] , \Z\R_DATA_TEMPR17[46] , 
        \Z\R_DATA_TEMPR18[46] , \Z\R_DATA_TEMPR19[46] , OR4_713_Y, 
        OR4_334_Y, OR4_114_Y, OR4_160_Y, OR4_287_Y, OR4_171_Y, 
        OR4_458_Y, OR4_704_Y, OR4_288_Y, OR4_585_Y, OR4_594_Y, 
        OR4_222_Y, OR2_29_Y, \Z\R_DATA_TEMPR22[18] , 
        \Z\R_DATA_TEMPR23[18] , OR4_649_Y, \Z\R_DATA_TEMPR12[19] , 
        \Z\R_DATA_TEMPR13[19] , \Z\R_DATA_TEMPR14[19] , 
        \Z\R_DATA_TEMPR15[19] , OR4_101_Y, \Z\R_DATA_TEMPR28[26] , 
        \Z\R_DATA_TEMPR29[26] , \Z\R_DATA_TEMPR30[26] , 
        \Z\R_DATA_TEMPR31[26] , OR4_589_Y, OR4_677_Y, OR4_480_Y, 
        OR4_384_Y, OR4_374_Y, OR4_569_Y, OR2_51_Y, 
        \Z\R_DATA_TEMPR22[24] , \Z\R_DATA_TEMPR23[24] , OR4_335_Y, 
        OR4_232_Y, OR4_376_Y, OR4_451_Y, OR4_270_Y, OR4_547_Y, 
        \Z\R_DATA_TEMPR28[34] , \Z\R_DATA_TEMPR29[34] , 
        \Z\R_DATA_TEMPR30[34] , \Z\R_DATA_TEMPR31[34] , OR4_117_Y, 
        OR4_195_Y, OR4_584_Y, OR4_137_Y, OR4_489_Y, 
        \Z\R_DATA_TEMPR20[60] , \Z\R_DATA_TEMPR20[61] , 
        \Z\R_DATA_TEMPR20[62] , \Z\R_DATA_TEMPR20[63] , 
        \Z\R_DATA_TEMPR20[64] , \Z\R_DATA_TEMPR20[65] , 
        \Z\R_DATA_TEMPR20[66] , \Z\R_DATA_TEMPR20[67] , 
        \Z\R_DATA_TEMPR20[68] , \Z\R_DATA_TEMPR20[69] , 
        \Z\R_DATA_TEMPR20[70] , \Z\R_DATA_TEMPR20[71] , 
        \Z\R_DATA_TEMPR20[72] , \Z\R_DATA_TEMPR20[73] , 
        \Z\R_DATA_TEMPR20[74] , \Z\R_DATA_TEMPR20[75] , 
        \Z\R_DATA_TEMPR20[76] , \Z\R_DATA_TEMPR20[77] , 
        \Z\R_DATA_TEMPR20[78] , \Z\R_DATA_TEMPR20[79] , 
        \Z\R_DATA_TEMPR20[41] , \Z\R_DATA_TEMPR20[42] , 
        \Z\R_DATA_TEMPR20[43] , \Z\R_DATA_TEMPR20[44] , 
        \Z\R_DATA_TEMPR20[45] , \Z\R_DATA_TEMPR20[46] , 
        \Z\R_DATA_TEMPR20[47] , \Z\R_DATA_TEMPR20[48] , 
        \Z\R_DATA_TEMPR20[49] , \Z\R_DATA_TEMPR20[50] , 
        \Z\R_DATA_TEMPR20[51] , \Z\R_DATA_TEMPR20[52] , 
        \Z\R_DATA_TEMPR20[53] , \Z\R_DATA_TEMPR20[54] , 
        \Z\R_DATA_TEMPR20[55] , \Z\R_DATA_TEMPR20[56] , 
        \Z\R_DATA_TEMPR20[57] , \Z\R_DATA_TEMPR20[58] , 
        \Z\R_DATA_TEMPR20[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C1_DB_DETECT, 
        \Z\ACCESS_BUSY[20][1] , OR4_304_Y, \Z\R_DATA_TEMPR4[59] , 
        \Z\R_DATA_TEMPR5[59] , \Z\R_DATA_TEMPR6[59] , 
        \Z\R_DATA_TEMPR7[59] , OR4_240_Y, OR4_347_Y, 
        \Z\R_DATA_TEMPR24[28] , \Z\R_DATA_TEMPR25[28] , 
        \Z\R_DATA_TEMPR26[28] , \Z\R_DATA_TEMPR27[28] , OR4_560_Y, 
        \Z\R_DATA_TEMPR28[9] , \Z\R_DATA_TEMPR29[9] , 
        \Z\R_DATA_TEMPR30[9] , \Z\R_DATA_TEMPR31[9] , OR4_63_Y, 
        \Z\R_DATA_TEMPR8[1] , \Z\R_DATA_TEMPR9[1] , 
        \Z\R_DATA_TEMPR11[1] , OR4_592_Y, \Z\R_DATA_TEMPR28[0] , 
        \Z\R_DATA_TEMPR29[0] , \Z\R_DATA_TEMPR30[0] , 
        \Z\R_DATA_TEMPR31[0] , OR4_168_Y, OR4_515_Y, OR4_27_Y, 
        OR4_118_Y, OR4_97_Y, \Z\R_DATA_TEMPR24[76] , 
        \Z\R_DATA_TEMPR25[76] , \Z\R_DATA_TEMPR26[76] , 
        \Z\R_DATA_TEMPR27[76] , \Z\R_DATA_TEMPR16[24] , 
        \Z\R_DATA_TEMPR17[24] , \Z\R_DATA_TEMPR18[24] , 
        \Z\R_DATA_TEMPR19[24] , OR4_46_Y, \Z\R_DATA_TEMPR16[47] , 
        \Z\R_DATA_TEMPR17[47] , \Z\R_DATA_TEMPR18[47] , 
        \Z\R_DATA_TEMPR19[47] , OR4_90_Y, OR4_239_Y, OR4_639_Y, 
        OR4_399_Y, OR4_157_Y, OR4_234_Y, OR4_667_Y, OR2_73_Y, 
        \Z\R_DATA_TEMPR22[75] , \Z\R_DATA_TEMPR23[75] , OR4_291_Y, 
        \Z\R_DATA_TEMPR8[45] , \Z\R_DATA_TEMPR9[45] , 
        \Z\R_DATA_TEMPR10[45] , \Z\R_DATA_TEMPR11[45] , OR2_18_Y, 
        \Z\R_DATA_TEMPR20[15] , \Z\R_DATA_TEMPR21[15] , OR4_468_Y, 
        OR4_198_Y, OR2_53_Y, \Z\R_DATA_TEMPR22[65] , 
        \Z\R_DATA_TEMPR23[65] , OR4_14_Y, \Z\R_DATA_TEMPR0[34] , 
        \Z\R_DATA_TEMPR1[34] , \Z\R_DATA_TEMPR2[34] , 
        \Z\R_DATA_TEMPR3[34] , \Z\R_DATA_TEMPR6[60] , 
        \Z\R_DATA_TEMPR6[61] , \Z\R_DATA_TEMPR6[62] , 
        \Z\R_DATA_TEMPR6[63] , \Z\R_DATA_TEMPR6[64] , 
        \Z\R_DATA_TEMPR6[65] , \Z\R_DATA_TEMPR6[66] , 
        \Z\R_DATA_TEMPR6[67] , \Z\R_DATA_TEMPR6[68] , 
        \Z\R_DATA_TEMPR6[69] , \Z\R_DATA_TEMPR6[70] , 
        \Z\R_DATA_TEMPR6[71] , \Z\R_DATA_TEMPR6[72] , 
        \Z\R_DATA_TEMPR6[73] , \Z\R_DATA_TEMPR6[74] , 
        \Z\R_DATA_TEMPR6[75] , \Z\R_DATA_TEMPR6[76] , 
        \Z\R_DATA_TEMPR6[77] , \Z\R_DATA_TEMPR6[78] , 
        \Z\R_DATA_TEMPR6[79] , \Z\R_DATA_TEMPR6[40] , 
        \Z\R_DATA_TEMPR6[41] , \Z\R_DATA_TEMPR6[42] , 
        \Z\R_DATA_TEMPR6[43] , \Z\R_DATA_TEMPR6[44] , 
        \Z\R_DATA_TEMPR6[45] , \Z\R_DATA_TEMPR6[46] , 
        \Z\R_DATA_TEMPR6[47] , \Z\R_DATA_TEMPR6[48] , 
        \Z\R_DATA_TEMPR6[49] , \Z\R_DATA_TEMPR6[50] , 
        \Z\R_DATA_TEMPR6[51] , \Z\R_DATA_TEMPR6[52] , 
        \Z\R_DATA_TEMPR6[53] , \Z\R_DATA_TEMPR6[54] , 
        \Z\R_DATA_TEMPR6[55] , \Z\R_DATA_TEMPR6[56] , 
        \Z\R_DATA_TEMPR6[57] , \Z\R_DATA_TEMPR6[58] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C1_DB_DETECT, 
        \Z\ACCESS_BUSY[6][1] , OR4_359_Y, \Z\R_DATA_TEMPR24[10] , 
        \Z\R_DATA_TEMPR25[10] , \Z\R_DATA_TEMPR26[10] , 
        \Z\R_DATA_TEMPR27[10] , OR4_461_Y, \Z\R_DATA_TEMPR16[52] , 
        \Z\R_DATA_TEMPR17[52] , \Z\R_DATA_TEMPR18[52] , 
        \Z\R_DATA_TEMPR19[52] , OR4_342_Y, \Z\R_DATA_TEMPR4[71] , 
        \Z\R_DATA_TEMPR5[71] , \Z\R_DATA_TEMPR7[71] , OR4_682_Y, 
        \Z\R_DATA_TEMPR24[17] , \Z\R_DATA_TEMPR25[17] , 
        \Z\R_DATA_TEMPR26[17] , \Z\R_DATA_TEMPR27[17] , OR2_78_Y, 
        \Z\R_DATA_TEMPR21[67] , \Z\R_DATA_TEMPR8[77] , 
        \Z\R_DATA_TEMPR9[77] , \Z\R_DATA_TEMPR10[77] , 
        \Z\R_DATA_TEMPR11[77] , \Z\R_DATA_TEMPR23[20] , 
        \Z\R_DATA_TEMPR23[22] , \Z\R_DATA_TEMPR23[23] , 
        \Z\R_DATA_TEMPR23[25] , \Z\R_DATA_TEMPR23[26] , 
        \Z\R_DATA_TEMPR23[27] , \Z\R_DATA_TEMPR23[28] , 
        \Z\R_DATA_TEMPR23[29] , \Z\R_DATA_TEMPR23[31] , 
        \Z\R_DATA_TEMPR23[32] , \Z\R_DATA_TEMPR23[33] , 
        \Z\R_DATA_TEMPR23[34] , \Z\R_DATA_TEMPR23[35] , 
        \Z\R_DATA_TEMPR23[36] , \Z\R_DATA_TEMPR23[37] , 
        \Z\R_DATA_TEMPR23[38] , \Z\R_DATA_TEMPR23[39] , 
        \Z\R_DATA_TEMPR23[0] , \Z\R_DATA_TEMPR23[1] , 
        \Z\R_DATA_TEMPR23[2] , \Z\R_DATA_TEMPR23[3] , 
        \Z\R_DATA_TEMPR23[4] , \Z\R_DATA_TEMPR23[5] , 
        \Z\R_DATA_TEMPR23[6] , \Z\R_DATA_TEMPR23[7] , 
        \Z\R_DATA_TEMPR23[8] , \Z\R_DATA_TEMPR23[9] , 
        \Z\R_DATA_TEMPR23[10] , \Z\R_DATA_TEMPR23[11] , 
        \Z\R_DATA_TEMPR23[12] , \Z\R_DATA_TEMPR23[13] , 
        \Z\R_DATA_TEMPR23[14] , \Z\R_DATA_TEMPR23[15] , 
        \Z\R_DATA_TEMPR23[16] , \Z\R_DATA_TEMPR23[17] , 
        \Z\R_DATA_TEMPR23[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0_DB_DETECT, 
        \Z\ACCESS_BUSY[23][0] , OR4_688_Y, OR4_105_Y, OR2_13_Y, 
        \Z\R_DATA_TEMPR22[5] , OR4_237_Y, \Z\R_DATA_TEMPR12[25] , 
        \Z\R_DATA_TEMPR13[25] , \Z\R_DATA_TEMPR14[25] , 
        \Z\R_DATA_TEMPR15[25] , OR4_676_Y, \Z\R_DATA_TEMPR8[36] , 
        \Z\R_DATA_TEMPR9[36] , \Z\R_DATA_TEMPR11[36] , OR4_716_Y, 
        OR2_41_Y, \Z\R_DATA_TEMPR22[62] , \Z\R_DATA_TEMPR23[62] , 
        OR4_161_Y, \Z\R_DATA_TEMPR0[75] , \Z\R_DATA_TEMPR1[75] , 
        \Z\R_DATA_TEMPR2[75] , \Z\R_DATA_TEMPR3[75] , OR4_446_Y, 
        \Z\R_DATA_TEMPR8[26] , \Z\R_DATA_TEMPR9[26] , 
        \Z\R_DATA_TEMPR11[26] , OR4_617_Y, \Z\R_DATA_TEMPR12[79] , 
        \Z\R_DATA_TEMPR13[79] , \Z\R_DATA_TEMPR14[79] , 
        \Z\R_DATA_TEMPR15[79] , OR4_715_Y, OR4_616_Y, 
        \Z\R_DATA_TEMPR22[67] , \Z\R_DATA_TEMPR23[67] , OR4_606_Y, 
        \Z\R_DATA_TEMPR16[69] , \Z\R_DATA_TEMPR17[69] , 
        \Z\R_DATA_TEMPR18[69] , \Z\R_DATA_TEMPR19[69] , OR4_364_Y, 
        \Z\R_DATA_TEMPR12[60] , \Z\R_DATA_TEMPR13[60] , 
        \Z\R_DATA_TEMPR14[60] , \Z\R_DATA_TEMPR15[60] , OR4_3_Y, 
        OR4_102_Y, OR2_72_Y, \Z\R_DATA_TEMPR22[70] , 
        \Z\R_DATA_TEMPR23[70] , OR4_54_Y, \Z\R_DATA_TEMPR28[70] , 
        \Z\R_DATA_TEMPR29[70] , \Z\R_DATA_TEMPR30[70] , 
        \Z\R_DATA_TEMPR31[70] , OR4_548_Y, \Z\R_DATA_TEMPR28[46] , 
        \Z\R_DATA_TEMPR29[46] , \Z\R_DATA_TEMPR30[46] , 
        \Z\R_DATA_TEMPR31[46] , OR4_96_Y, \Z\R_DATA_TEMPR4[7] , 
        \Z\R_DATA_TEMPR6[7] , \Z\R_DATA_TEMPR7[7] , OR4_283_Y, 
        \Z\R_DATA_TEMPR24[64] , \Z\R_DATA_TEMPR25[64] , 
        \Z\R_DATA_TEMPR26[64] , \Z\R_DATA_TEMPR27[64] , OR4_571_Y, 
        OR4_205_Y, OR4_472_Y, OR4_274_Y, OR4_450_Y, 
        \Z\R_DATA_TEMPR12[27] , \Z\R_DATA_TEMPR13[27] , 
        \Z\R_DATA_TEMPR14[27] , \Z\R_DATA_TEMPR15[27] , OR4_611_Y, 
        OR4_419_Y, OR4_366_Y, OR2_28_Y, \Z\R_DATA_TEMPR20[14] , 
        \Z\R_DATA_TEMPR21[14] , OR4_351_Y, \Z\R_DATA_TEMPR4[70] , 
        \Z\R_DATA_TEMPR5[70] , \Z\R_DATA_TEMPR7[70] , OR4_624_Y, 
        \Z\R_DATA_TEMPR24[27] , \Z\R_DATA_TEMPR25[27] , 
        \Z\R_DATA_TEMPR26[27] , \Z\R_DATA_TEMPR27[27] , OR4_637_Y, 
        \Z\R_DATA_TEMPR16[25] , \Z\R_DATA_TEMPR17[25] , 
        \Z\R_DATA_TEMPR18[25] , \Z\R_DATA_TEMPR19[25] , OR4_72_Y, 
        \Z\R_DATA_TEMPR0[50] , \Z\R_DATA_TEMPR1[50] , 
        \Z\R_DATA_TEMPR2[50] , \Z\R_DATA_TEMPR3[50] , OR4_119_Y, 
        \Z\R_DATA_TEMPR24[37] , \Z\R_DATA_TEMPR25[37] , 
        \Z\R_DATA_TEMPR26[37] , \Z\R_DATA_TEMPR27[37] , OR4_226_Y, 
        \Z\R_DATA_TEMPR4[64] , \Z\R_DATA_TEMPR5[64] , 
        \Z\R_DATA_TEMPR7[64] , OR4_546_Y, \Z\R_DATA_TEMPR28[65] , 
        \Z\R_DATA_TEMPR29[65] , \Z\R_DATA_TEMPR30[65] , 
        \Z\R_DATA_TEMPR31[65] , OR4_554_Y, \Z\R_DATA_TEMPR4[27] , 
        \Z\R_DATA_TEMPR6[27] , \Z\R_DATA_TEMPR7[27] , OR4_629_Y, 
        \Z\R_DATA_TEMPR0[26] , \Z\R_DATA_TEMPR1[26] , 
        \Z\R_DATA_TEMPR2[26] , \Z\R_DATA_TEMPR3[26] , 
        \Z\R_DATA_TEMPR4[24] , \Z\R_DATA_TEMPR6[24] , 
        \Z\R_DATA_TEMPR7[24] , OR2_17_Y, \Z\R_DATA_TEMPR21[55] , 
        OR4_178_Y, OR4_373_Y, OR4_314_Y, OR4_371_Y, OR4_181_Y, 
        OR4_520_Y, OR4_70_Y, OR4_597_Y, OR2_10_Y, 
        \Z\R_DATA_TEMPR20[9] , \Z\R_DATA_TEMPR21[9] , OR4_318_Y, 
        \Z\R_DATA_TEMPR8[79] , \Z\R_DATA_TEMPR9[79] , 
        \Z\R_DATA_TEMPR10[79] , \Z\R_DATA_TEMPR11[79] , OR4_527_Y, 
        \Z\R_DATA_TEMPR4[32] , \Z\R_DATA_TEMPR6[32] , 
        \Z\R_DATA_TEMPR7[32] , OR4_672_Y, OR4_360_Y, OR2_14_Y, 
        \Z\R_DATA_TEMPR22[32] , OR4_220_Y, \Z\R_DATA_TEMPR12[78] , 
        \Z\R_DATA_TEMPR13[78] , \Z\R_DATA_TEMPR14[78] , 
        \Z\R_DATA_TEMPR15[78] , OR2_77_Y, \Z\R_DATA_TEMPR21[42] , 
        OR4_552_Y, \Z\R_DATA_TEMPR4[25] , \Z\R_DATA_TEMPR6[25] , 
        \Z\R_DATA_TEMPR7[25] , OR4_690_Y, OR4_567_Y, OR4_255_Y, 
        OR4_602_Y, \Z\R_DATA_TEMPR16[74] , \Z\R_DATA_TEMPR17[74] , 
        \Z\R_DATA_TEMPR18[74] , \Z\R_DATA_TEMPR19[74] , OR4_678_Y, 
        \Z\R_DATA_TEMPR12[37] , \Z\R_DATA_TEMPR13[37] , 
        \Z\R_DATA_TEMPR14[37] , \Z\R_DATA_TEMPR15[37] , OR2_70_Y, 
        \Z\R_DATA_TEMPR21[43] , OR4_694_Y, \Z\R_DATA_TEMPR4[48] , 
        \Z\R_DATA_TEMPR5[48] , \Z\R_DATA_TEMPR7[48] , 
        \Z\R_DATA_TEMPR18[21] , \Z\R_DATA_TEMPR18[22] , 
        \Z\R_DATA_TEMPR18[23] , \Z\R_DATA_TEMPR18[26] , 
        \Z\R_DATA_TEMPR18[27] , \Z\R_DATA_TEMPR18[28] , 
        \Z\R_DATA_TEMPR18[29] , \Z\R_DATA_TEMPR18[30] , 
        \Z\R_DATA_TEMPR18[31] , \Z\R_DATA_TEMPR18[32] , 
        \Z\R_DATA_TEMPR18[33] , \Z\R_DATA_TEMPR18[34] , 
        \Z\R_DATA_TEMPR18[36] , \Z\R_DATA_TEMPR18[37] , 
        \Z\R_DATA_TEMPR18[38] , \Z\R_DATA_TEMPR18[39] , 
        \Z\R_DATA_TEMPR18[0] , \Z\R_DATA_TEMPR18[1] , 
        \Z\R_DATA_TEMPR18[3] , \Z\R_DATA_TEMPR18[4] , 
        \Z\R_DATA_TEMPR18[5] , \Z\R_DATA_TEMPR18[6] , 
        \Z\R_DATA_TEMPR18[7] , \Z\R_DATA_TEMPR18[8] , 
        \Z\R_DATA_TEMPR18[9] , \Z\R_DATA_TEMPR18[10] , 
        \Z\R_DATA_TEMPR18[11] , \Z\R_DATA_TEMPR18[12] , 
        \Z\R_DATA_TEMPR18[13] , \Z\R_DATA_TEMPR18[14] , 
        \Z\R_DATA_TEMPR18[15] , \Z\R_DATA_TEMPR18[16] , 
        \Z\R_DATA_TEMPR18[17] , \Z\R_DATA_TEMPR18[18] , 
        \Z\R_DATA_TEMPR18[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0_DB_DETECT, 
        \Z\ACCESS_BUSY[18][0] , OR4_144_Y, \Z\R_DATA_TEMPR12[12] , 
        \Z\R_DATA_TEMPR13[12] , \Z\R_DATA_TEMPR14[12] , 
        \Z\R_DATA_TEMPR15[12] , OR4_608_Y, OR4_245_Y, OR4_17_Y, 
        OR4_52_Y, OR4_192_Y, OR4_116_Y, \Z\R_DATA_TEMPR0[33] , 
        \Z\R_DATA_TEMPR1[33] , \Z\R_DATA_TEMPR2[33] , 
        \Z\R_DATA_TEMPR3[33] , \Z\R_DATA_TEMPR14[61] , 
        \Z\R_DATA_TEMPR14[63] , \Z\R_DATA_TEMPR14[64] , 
        \Z\R_DATA_TEMPR14[65] , \Z\R_DATA_TEMPR14[66] , 
        \Z\R_DATA_TEMPR14[67] , \Z\R_DATA_TEMPR14[68] , 
        \Z\R_DATA_TEMPR14[69] , \Z\R_DATA_TEMPR14[70] , 
        \Z\R_DATA_TEMPR14[71] , \Z\R_DATA_TEMPR14[72] , 
        \Z\R_DATA_TEMPR14[73] , \Z\R_DATA_TEMPR14[74] , 
        \Z\R_DATA_TEMPR14[75] , \Z\R_DATA_TEMPR14[76] , 
        \Z\R_DATA_TEMPR14[77] , \Z\R_DATA_TEMPR14[40] , 
        \Z\R_DATA_TEMPR14[41] , \Z\R_DATA_TEMPR14[43] , 
        \Z\R_DATA_TEMPR14[44] , \Z\R_DATA_TEMPR14[45] , 
        \Z\R_DATA_TEMPR14[46] , \Z\R_DATA_TEMPR14[47] , 
        \Z\R_DATA_TEMPR14[48] , \Z\R_DATA_TEMPR14[49] , 
        \Z\R_DATA_TEMPR14[50] , \Z\R_DATA_TEMPR14[51] , 
        \Z\R_DATA_TEMPR14[52] , \Z\R_DATA_TEMPR14[53] , 
        \Z\R_DATA_TEMPR14[54] , \Z\R_DATA_TEMPR14[55] , 
        \Z\R_DATA_TEMPR14[56] , \Z\R_DATA_TEMPR14[57] , 
        \Z\R_DATA_TEMPR14[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C1_DB_DETECT, 
        \Z\ACCESS_BUSY[14][1] , OR4_139_Y, \Z\R_DATA_TEMPR28[23] , 
        \Z\R_DATA_TEMPR29[23] , \Z\R_DATA_TEMPR30[23] , 
        \Z\R_DATA_TEMPR31[23] , OR4_79_Y, \Z\R_DATA_TEMPR8[50] , 
        \Z\R_DATA_TEMPR9[50] , \Z\R_DATA_TEMPR10[50] , 
        \Z\R_DATA_TEMPR11[50] , \Z\R_DATA_TEMPR11[20] , 
        \Z\R_DATA_TEMPR11[21] , \Z\R_DATA_TEMPR11[22] , 
        \Z\R_DATA_TEMPR11[23] , \Z\R_DATA_TEMPR11[24] , 
        \Z\R_DATA_TEMPR11[25] , \Z\R_DATA_TEMPR11[28] , 
        \Z\R_DATA_TEMPR11[29] , \Z\R_DATA_TEMPR11[30] , 
        \Z\R_DATA_TEMPR11[31] , \Z\R_DATA_TEMPR11[32] , 
        \Z\R_DATA_TEMPR11[33] , \Z\R_DATA_TEMPR11[34] , 
        \Z\R_DATA_TEMPR11[35] , \Z\R_DATA_TEMPR11[37] , 
        \Z\R_DATA_TEMPR11[38] , \Z\R_DATA_TEMPR11[39] , 
        \Z\R_DATA_TEMPR11[0] , \Z\R_DATA_TEMPR11[3] , 
        \Z\R_DATA_TEMPR11[4] , \Z\R_DATA_TEMPR11[5] , 
        \Z\R_DATA_TEMPR11[6] , \Z\R_DATA_TEMPR11[7] , 
        \Z\R_DATA_TEMPR11[8] , \Z\R_DATA_TEMPR11[9] , 
        \Z\R_DATA_TEMPR11[10] , \Z\R_DATA_TEMPR11[11] , 
        \Z\R_DATA_TEMPR11[12] , \Z\R_DATA_TEMPR11[13] , 
        \Z\R_DATA_TEMPR11[14] , \Z\R_DATA_TEMPR11[15] , 
        \Z\R_DATA_TEMPR11[17] , \Z\R_DATA_TEMPR11[18] , 
        \Z\R_DATA_TEMPR11[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0_DB_DETECT, 
        \Z\ACCESS_BUSY[11][0] , OR4_251_Y, \Z\R_DATA_TEMPR16[55] , 
        \Z\R_DATA_TEMPR17[55] , \Z\R_DATA_TEMPR18[55] , 
        \Z\R_DATA_TEMPR19[55] , OR4_285_Y, OR2_6_Y, 
        \Z\R_DATA_TEMPR22[33] , OR4_296_Y, \Z\R_DATA_TEMPR12[49] , 
        \Z\R_DATA_TEMPR13[49] , \Z\R_DATA_TEMPR15[49] , OR4_412_Y, 
        OR4_654_Y, OR4_507_Y, OR4_498_Y, OR4_227_Y, OR4_583_Y, 
        \Z\R_DATA_TEMPR4[75] , \Z\R_DATA_TEMPR5[75] , 
        \Z\R_DATA_TEMPR7[75] , OR4_12_Y, \Z\R_DATA_TEMPR0[58] , 
        \Z\R_DATA_TEMPR1[58] , \Z\R_DATA_TEMPR2[58] , 
        \Z\R_DATA_TEMPR3[58] , \Z\R_DATA_TEMPR19[21] , 
        \Z\R_DATA_TEMPR19[22] , \Z\R_DATA_TEMPR19[23] , 
        \Z\R_DATA_TEMPR19[26] , \Z\R_DATA_TEMPR19[27] , 
        \Z\R_DATA_TEMPR19[28] , \Z\R_DATA_TEMPR19[29] , 
        \Z\R_DATA_TEMPR19[30] , \Z\R_DATA_TEMPR19[31] , 
        \Z\R_DATA_TEMPR19[32] , \Z\R_DATA_TEMPR19[33] , 
        \Z\R_DATA_TEMPR19[34] , \Z\R_DATA_TEMPR19[36] , 
        \Z\R_DATA_TEMPR19[37] , \Z\R_DATA_TEMPR19[38] , 
        \Z\R_DATA_TEMPR19[39] , \Z\R_DATA_TEMPR19[0] , 
        \Z\R_DATA_TEMPR19[1] , \Z\R_DATA_TEMPR19[3] , 
        \Z\R_DATA_TEMPR19[4] , \Z\R_DATA_TEMPR19[5] , 
        \Z\R_DATA_TEMPR19[6] , \Z\R_DATA_TEMPR19[7] , 
        \Z\R_DATA_TEMPR19[8] , \Z\R_DATA_TEMPR19[9] , 
        \Z\R_DATA_TEMPR19[10] , \Z\R_DATA_TEMPR19[11] , 
        \Z\R_DATA_TEMPR19[12] , \Z\R_DATA_TEMPR19[13] , 
        \Z\R_DATA_TEMPR19[14] , \Z\R_DATA_TEMPR19[15] , 
        \Z\R_DATA_TEMPR19[16] , \Z\R_DATA_TEMPR19[17] , 
        \Z\R_DATA_TEMPR19[18] , \Z\R_DATA_TEMPR19[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0_DB_DETECT, 
        \Z\ACCESS_BUSY[19][0] , OR4_699_Y, \Z\R_DATA_TEMPR4[74] , 
        \Z\R_DATA_TEMPR5[74] , \Z\R_DATA_TEMPR7[74] , OR4_710_Y, 
        \Z\R_DATA_TEMPR12[61] , \Z\R_DATA_TEMPR13[61] , 
        \Z\R_DATA_TEMPR15[61] , OR4_322_Y, \Z\R_DATA_TEMPR4[72] , 
        \Z\R_DATA_TEMPR5[72] , \Z\R_DATA_TEMPR7[72] , OR4_313_Y, 
        \Z\R_DATA_TEMPR4[18] , \Z\R_DATA_TEMPR6[18] , 
        \Z\R_DATA_TEMPR7[18] , OR4_473_Y, OR4_657_Y, OR4_717_Y, 
        OR4_273_Y, \Z\R_DATA_TEMPR4[47] , \Z\R_DATA_TEMPR5[47] , 
        \Z\R_DATA_TEMPR7[47] , OR4_338_Y, OR4_111_Y, OR4_574_Y, 
        OR4_609_Y, \Z\R_DATA_TEMPR28[55] , \Z\R_DATA_TEMPR29[55] , 
        \Z\R_DATA_TEMPR30[55] , \Z\R_DATA_TEMPR31[55] , OR4_290_Y, 
        \Z\R_DATA_TEMPR24[59] , \Z\R_DATA_TEMPR25[59] , 
        \Z\R_DATA_TEMPR26[59] , \Z\R_DATA_TEMPR27[59] , OR4_203_Y, 
        \Z\R_DATA_TEMPR12[59] , \Z\R_DATA_TEMPR13[59] , 
        \Z\R_DATA_TEMPR15[59] , \Z\R_DATA_TEMPR9[20] , 
        \Z\R_DATA_TEMPR9[21] , \Z\R_DATA_TEMPR9[22] , 
        \Z\R_DATA_TEMPR9[23] , \Z\R_DATA_TEMPR9[24] , 
        \Z\R_DATA_TEMPR9[25] , \Z\R_DATA_TEMPR9[28] , 
        \Z\R_DATA_TEMPR9[29] , \Z\R_DATA_TEMPR9[30] , 
        \Z\R_DATA_TEMPR9[31] , \Z\R_DATA_TEMPR9[32] , 
        \Z\R_DATA_TEMPR9[33] , \Z\R_DATA_TEMPR9[34] , 
        \Z\R_DATA_TEMPR9[35] , \Z\R_DATA_TEMPR9[37] , 
        \Z\R_DATA_TEMPR9[38] , \Z\R_DATA_TEMPR9[39] , 
        \Z\R_DATA_TEMPR9[0] , \Z\R_DATA_TEMPR9[3] , 
        \Z\R_DATA_TEMPR9[4] , \Z\R_DATA_TEMPR9[5] , 
        \Z\R_DATA_TEMPR9[6] , \Z\R_DATA_TEMPR9[7] , 
        \Z\R_DATA_TEMPR9[8] , \Z\R_DATA_TEMPR9[9] , 
        \Z\R_DATA_TEMPR9[10] , \Z\R_DATA_TEMPR9[11] , 
        \Z\R_DATA_TEMPR9[12] , \Z\R_DATA_TEMPR9[13] , 
        \Z\R_DATA_TEMPR9[14] , \Z\R_DATA_TEMPR9[15] , 
        \Z\R_DATA_TEMPR9[17] , \Z\R_DATA_TEMPR9[18] , 
        \Z\R_DATA_TEMPR9[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0_DB_DETECT, 
        \Z\ACCESS_BUSY[9][0] , OR4_426_Y, \Z\R_DATA_TEMPR0[67] , 
        \Z\R_DATA_TEMPR1[67] , \Z\R_DATA_TEMPR2[67] , 
        \Z\R_DATA_TEMPR3[67] , OR2_27_Y, \Z\R_DATA_TEMPR21[58] , 
        OR2_16_Y, \Z\R_DATA_TEMPR21[48] , OR2_20_Y, 
        \Z\R_DATA_TEMPR21[66] , OR4_136_Y, OR4_56_Y, OR2_62_Y, 
        \Z\R_DATA_TEMPR22[4] , OR4_346_Y, \Z\R_DATA_TEMPR8[54] , 
        \Z\R_DATA_TEMPR9[54] , \Z\R_DATA_TEMPR10[54] , 
        \Z\R_DATA_TEMPR11[54] , OR4_439_Y, OR4_15_Y, OR4_267_Y, 
        OR4_566_Y, OR4_134_Y, OR4_662_Y, OR4_432_Y, OR4_289_Y, 
        \Z\R_DATA_TEMPR8[56] , \Z\R_DATA_TEMPR9[56] , 
        \Z\R_DATA_TEMPR10[56] , \Z\R_DATA_TEMPR11[56] , OR2_76_Y, 
        \Z\R_DATA_TEMPR20[13] , \Z\R_DATA_TEMPR21[13] , OR4_528_Y, 
        \Z\R_DATA_TEMPR8[13] , \Z\R_DATA_TEMPR0[78] , 
        \Z\R_DATA_TEMPR1[78] , \Z\R_DATA_TEMPR2[78] , 
        \Z\R_DATA_TEMPR3[78] , OR4_444_Y, \Z\R_DATA_TEMPR12[68] , 
        \Z\R_DATA_TEMPR13[68] , \Z\R_DATA_TEMPR15[68] , OR4_510_Y, 
        \Z\R_DATA_TEMPR24[46] , \Z\R_DATA_TEMPR25[46] , 
        \Z\R_DATA_TEMPR26[46] , \Z\R_DATA_TEMPR27[46] , OR4_668_Y, 
        \Z\R_DATA_TEMPR16[57] , \Z\R_DATA_TEMPR17[57] , 
        \Z\R_DATA_TEMPR18[57] , \Z\R_DATA_TEMPR19[57] , 
        \Z\R_DATA_TEMPR17[60] , \Z\R_DATA_TEMPR17[61] , 
        \Z\R_DATA_TEMPR17[63] , \Z\R_DATA_TEMPR17[64] , 
        \Z\R_DATA_TEMPR17[65] , \Z\R_DATA_TEMPR17[66] , 
        \Z\R_DATA_TEMPR17[67] , \Z\R_DATA_TEMPR17[68] , 
        \Z\R_DATA_TEMPR17[70] , \Z\R_DATA_TEMPR17[71] , 
        \Z\R_DATA_TEMPR17[72] , \Z\R_DATA_TEMPR17[73] , 
        \Z\R_DATA_TEMPR17[75] , \Z\R_DATA_TEMPR17[76] , 
        \Z\R_DATA_TEMPR17[77] , \Z\R_DATA_TEMPR17[78] , 
        \Z\R_DATA_TEMPR17[79] , \Z\R_DATA_TEMPR17[40] , 
        \Z\R_DATA_TEMPR17[41] , \Z\R_DATA_TEMPR17[43] , 
        \Z\R_DATA_TEMPR17[44] , \Z\R_DATA_TEMPR17[45] , 
        \Z\R_DATA_TEMPR17[48] , \Z\R_DATA_TEMPR17[49] , 
        \Z\R_DATA_TEMPR17[50] , \Z\R_DATA_TEMPR17[51] , 
        \Z\R_DATA_TEMPR17[53] , \Z\R_DATA_TEMPR17[54] , 
        \Z\R_DATA_TEMPR17[56] , \Z\R_DATA_TEMPR17[58] , 
        \Z\R_DATA_TEMPR17[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C1_DB_DETECT, 
        \Z\ACCESS_BUSY[17][1] , OR4_519_Y, \Z\R_DATA_TEMPR8[39] , 
        \Z\R_DATA_TEMPR16[63] , \Z\R_DATA_TEMPR18[63] , 
        \Z\R_DATA_TEMPR19[63] , OR4_41_Y, \Z\R_DATA_TEMPR16[49] , 
        \Z\R_DATA_TEMPR18[49] , \Z\R_DATA_TEMPR19[49] , OR4_19_Y, 
        OR4_147_Y, OR4_576_Y, OR4_0_Y, OR4_392_Y, OR4_474_Y, OR4_231_Y, 
        OR4_215_Y, OR4_389_Y, \Z\R_DATA_TEMPR16[53] , 
        \Z\R_DATA_TEMPR18[53] , \Z\R_DATA_TEMPR19[53] , OR4_599_Y, 
        OR4_680_Y, OR4_452_Y, OR4_418_Y, OR2_30_Y, 
        \Z\R_DATA_TEMPR22[35] , OR4_496_Y, \Z\R_DATA_TEMPR16[43] , 
        \Z\R_DATA_TEMPR18[43] , \Z\R_DATA_TEMPR19[43] , OR4_411_Y, 
        \Z\R_DATA_TEMPR12[52] , \Z\R_DATA_TEMPR13[52] , 
        \Z\R_DATA_TEMPR15[52] , \Z\R_DATA_TEMPR8[22] , OR4_526_Y, 
        OR4_656_Y, OR4_356_Y, OR4_508_Y, OR4_263_Y, OR4_355_Y, 
        OR2_50_Y, \Z\R_DATA_TEMPR22[60] , \Z\R_DATA_TEMPR23[60] , 
        OR4_530_Y, OR4_591_Y, OR4_545_Y, OR4_162_Y, OR4_59_Y, 
        \Z\R_DATA_TEMPR0[64] , \Z\R_DATA_TEMPR1[64] , 
        \Z\R_DATA_TEMPR2[64] , \Z\R_DATA_TEMPR3[64] , 
        \Z\R_DATA_TEMPR16[60] , \Z\R_DATA_TEMPR16[61] , 
        \Z\R_DATA_TEMPR16[64] , \Z\R_DATA_TEMPR16[65] , 
        \Z\R_DATA_TEMPR16[66] , \Z\R_DATA_TEMPR16[67] , 
        \Z\R_DATA_TEMPR16[68] , \Z\R_DATA_TEMPR16[70] , 
        \Z\R_DATA_TEMPR16[71] , \Z\R_DATA_TEMPR16[72] , 
        \Z\R_DATA_TEMPR16[73] , \Z\R_DATA_TEMPR16[75] , 
        \Z\R_DATA_TEMPR16[76] , \Z\R_DATA_TEMPR16[77] , 
        \Z\R_DATA_TEMPR16[78] , \Z\R_DATA_TEMPR16[79] , 
        \Z\R_DATA_TEMPR16[40] , \Z\R_DATA_TEMPR16[41] , 
        \Z\R_DATA_TEMPR16[44] , \Z\R_DATA_TEMPR16[45] , 
        \Z\R_DATA_TEMPR16[48] , \Z\R_DATA_TEMPR16[50] , 
        \Z\R_DATA_TEMPR16[51] , \Z\R_DATA_TEMPR16[54] , 
        \Z\R_DATA_TEMPR16[56] , \Z\R_DATA_TEMPR16[58] , 
        \Z\R_DATA_TEMPR16[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C1_DB_DETECT, 
        \Z\ACCESS_BUSY[16][1] , OR4_598_Y, \Z\R_DATA_TEMPR28[64] , 
        \Z\R_DATA_TEMPR29[64] , \Z\R_DATA_TEMPR30[64] , 
        \Z\R_DATA_TEMPR31[64] , \Z\R_DATA_TEMPR0[48] , 
        \Z\R_DATA_TEMPR1[48] , \Z\R_DATA_TEMPR2[48] , 
        \Z\R_DATA_TEMPR3[48] , OR2_26_Y, \Z\R_DATA_TEMPR21[54] , 
        OR4_539_Y, \Z\R_DATA_TEMPR0[10] , \Z\R_DATA_TEMPR1[10] , 
        \Z\R_DATA_TEMPR2[10] , \Z\R_DATA_TEMPR3[10] , OR4_573_Y, 
        \Z\R_DATA_TEMPR0[0] , \Z\R_DATA_TEMPR1[0] , 
        \Z\R_DATA_TEMPR2[0] , \Z\R_DATA_TEMPR3[0] , OR4_43_Y, OR2_45_Y, 
        \Z\R_DATA_TEMPR22[57] , \Z\R_DATA_TEMPR23[57] , 
        \Z\R_DATA_TEMPR20[20] , \Z\R_DATA_TEMPR20[21] , 
        \Z\R_DATA_TEMPR20[22] , \Z\R_DATA_TEMPR20[23] , 
        \Z\R_DATA_TEMPR20[24] , \Z\R_DATA_TEMPR20[25] , 
        \Z\R_DATA_TEMPR20[26] , \Z\R_DATA_TEMPR20[27] , 
        \Z\R_DATA_TEMPR20[28] , \Z\R_DATA_TEMPR20[29] , 
        \Z\R_DATA_TEMPR20[31] , \Z\R_DATA_TEMPR20[32] , 
        \Z\R_DATA_TEMPR20[33] , \Z\R_DATA_TEMPR20[34] , 
        \Z\R_DATA_TEMPR20[35] , \Z\R_DATA_TEMPR20[36] , 
        \Z\R_DATA_TEMPR20[37] , \Z\R_DATA_TEMPR20[38] , 
        \Z\R_DATA_TEMPR20[39] , \Z\R_DATA_TEMPR20[0] , 
        \Z\R_DATA_TEMPR20[1] , \Z\R_DATA_TEMPR20[2] , 
        \Z\R_DATA_TEMPR20[3] , \Z\R_DATA_TEMPR20[4] , 
        \Z\R_DATA_TEMPR20[5] , \Z\R_DATA_TEMPR20[6] , 
        \Z\R_DATA_TEMPR20[7] , \Z\R_DATA_TEMPR20[8] , 
        \Z\R_DATA_TEMPR20[10] , \Z\R_DATA_TEMPR20[11] , 
        \Z\R_DATA_TEMPR20[12] , \Z\R_DATA_TEMPR20[16] , 
        \Z\R_DATA_TEMPR20[17] , \Z\R_DATA_TEMPR20[18] , 
        \Z\R_DATA_TEMPR20[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0_DB_DETECT, 
        \Z\ACCESS_BUSY[20][0] , \Z\R_DATA_TEMPR24[3] , 
        \Z\R_DATA_TEMPR25[3] , \Z\R_DATA_TEMPR26[3] , 
        \Z\R_DATA_TEMPR27[3] , OR4_503_Y, \Z\R_DATA_TEMPR12[65] , 
        \Z\R_DATA_TEMPR13[65] , \Z\R_DATA_TEMPR15[65] , 
        \Z\R_DATA_TEMPR24[1] , \Z\R_DATA_TEMPR25[1] , 
        \Z\R_DATA_TEMPR26[1] , \Z\R_DATA_TEMPR27[1] , OR4_309_Y, 
        OR4_705_Y, OR4_141_Y, \Z\R_DATA_TEMPR0[73] , 
        \Z\R_DATA_TEMPR1[73] , \Z\R_DATA_TEMPR2[73] , 
        \Z\R_DATA_TEMPR3[73] , OR2_3_Y, \Z\R_DATA_TEMPR21[71] , 
        OR4_381_Y, OR2_59_Y, \Z\R_DATA_TEMPR22[46] , 
        \Z\R_DATA_TEMPR23[46] , OR4_709_Y, \Z\R_DATA_TEMPR4[33] , 
        \Z\R_DATA_TEMPR6[33] , \Z\R_DATA_TEMPR7[33] , OR4_438_Y, 
        \Z\R_DATA_TEMPR4[76] , \Z\R_DATA_TEMPR5[76] , 
        \Z\R_DATA_TEMPR7[76] , OR4_124_Y, \Z\R_DATA_TEMPR12[66] , 
        \Z\R_DATA_TEMPR13[66] , \Z\R_DATA_TEMPR15[66] , OR4_91_Y, 
        \Z\R_DATA_TEMPR0[32] , \Z\R_DATA_TEMPR1[32] , 
        \Z\R_DATA_TEMPR2[32] , \Z\R_DATA_TEMPR3[32] , OR4_562_Y, 
        OR4_323_Y, OR4_431_Y, \Z\R_DATA_TEMPR28[56] , 
        \Z\R_DATA_TEMPR29[56] , \Z\R_DATA_TEMPR30[56] , 
        \Z\R_DATA_TEMPR31[56] , \Z\R_DATA_TEMPR21[33] , 
        \Z\R_DATA_TEMPR4[53] , \Z\R_DATA_TEMPR5[53] , 
        \Z\R_DATA_TEMPR7[53] , OR2_0_Y, \Z\R_DATA_TEMPR21[74] , 
        OR4_256_Y, OR4_199_Y, OR4_35_Y, OR4_207_Y, OR4_523_Y, 
        OR4_393_Y, OR4_252_Y, OR4_202_Y, OR4_58_Y, 
        \Z\R_DATA_TEMPR0[22] , \Z\R_DATA_TEMPR1[22] , 
        \Z\R_DATA_TEMPR2[22] , \Z\R_DATA_TEMPR3[22] , OR4_659_Y, 
        \Z\R_DATA_TEMPR0[76] , \Z\R_DATA_TEMPR1[76] , 
        \Z\R_DATA_TEMPR2[76] , \Z\R_DATA_TEMPR3[76] , 
        \Z\R_DATA_TEMPR4[77] , \Z\R_DATA_TEMPR5[77] , 
        \Z\R_DATA_TEMPR7[77] , OR4_131_Y, OR4_651_Y, OR4_414_Y, 
        \Z\R_DATA_TEMPR18[60] , \Z\R_DATA_TEMPR18[61] , 
        \Z\R_DATA_TEMPR18[64] , \Z\R_DATA_TEMPR18[65] , 
        \Z\R_DATA_TEMPR18[66] , \Z\R_DATA_TEMPR18[67] , 
        \Z\R_DATA_TEMPR18[68] , \Z\R_DATA_TEMPR18[70] , 
        \Z\R_DATA_TEMPR18[71] , \Z\R_DATA_TEMPR18[72] , 
        \Z\R_DATA_TEMPR18[73] , \Z\R_DATA_TEMPR18[75] , 
        \Z\R_DATA_TEMPR18[76] , \Z\R_DATA_TEMPR18[77] , 
        \Z\R_DATA_TEMPR18[78] , \Z\R_DATA_TEMPR18[79] , 
        \Z\R_DATA_TEMPR18[40] , \Z\R_DATA_TEMPR18[41] , 
        \Z\R_DATA_TEMPR18[44] , \Z\R_DATA_TEMPR18[45] , 
        \Z\R_DATA_TEMPR18[48] , \Z\R_DATA_TEMPR18[50] , 
        \Z\R_DATA_TEMPR18[51] , \Z\R_DATA_TEMPR18[54] , 
        \Z\R_DATA_TEMPR18[56] , \Z\R_DATA_TEMPR18[58] , 
        \Z\R_DATA_TEMPR18[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C1_DB_DETECT, 
        \Z\ACCESS_BUSY[18][1] , OR4_700_Y, OR4_664_Y, OR4_674_Y, 
        OR4_447_Y, \Z\R_DATA_TEMPR0[46] , \Z\R_DATA_TEMPR1[46] , 
        \Z\R_DATA_TEMPR2[46] , \Z\R_DATA_TEMPR3[46] , OR2_4_Y, 
        \Z\R_DATA_TEMPR21[12] , OR4_557_Y, \Z\R_DATA_TEMPR12[55] , 
        \Z\R_DATA_TEMPR13[55] , \Z\R_DATA_TEMPR15[55] , OR4_250_Y, 
        OR4_442_Y, OR2_31_Y, \Z\R_DATA_TEMPR22[51] , 
        \Z\R_DATA_TEMPR23[51] , OR4_379_Y, \Z\R_DATA_TEMPR0[37] , 
        \Z\R_DATA_TEMPR1[37] , \Z\R_DATA_TEMPR2[37] , 
        \Z\R_DATA_TEMPR3[37] , OR4_8_Y, \Z\R_DATA_TEMPR4[42] , 
        \Z\R_DATA_TEMPR5[42] , \Z\R_DATA_TEMPR7[42] , OR4_24_Y, 
        \Z\R_DATA_TEMPR24[19] , \Z\R_DATA_TEMPR25[19] , 
        \Z\R_DATA_TEMPR26[19] , \Z\R_DATA_TEMPR27[19] , OR4_582_Y, 
        \Z\R_DATA_TEMPR8[25] , OR4_487_Y, OR4_613_Y, 
        \Z\R_DATA_TEMPR19[67] , OR4_93_Y, \Z\R_DATA_TEMPR12[64] , 
        \Z\R_DATA_TEMPR13[64] , \Z\R_DATA_TEMPR15[64] , OR4_563_Y, 
        \Z\R_DATA_TEMPR16[37] , \Z\R_DATA_TEMPR17[37] , OR4_326_Y, 
        \Z\R_DATA_TEMPR28[78] , \Z\R_DATA_TEMPR29[78] , 
        \Z\R_DATA_TEMPR30[78] , \Z\R_DATA_TEMPR31[78] , OR4_369_Y, 
        OR4_186_Y, OR4_257_Y, OR4_194_Y, \Z\R_DATA_TEMPR24[45] , 
        \Z\R_DATA_TEMPR25[45] , \Z\R_DATA_TEMPR26[45] , 
        \Z\R_DATA_TEMPR27[45] , OR4_281_Y, \Z\R_DATA_TEMPR19[44] , 
        OR4_424_Y, \Z\R_DATA_TEMPR19[68] , \Z\R_DATA_TEMPR0[69] , 
        \Z\R_DATA_TEMPR1[69] , \Z\R_DATA_TEMPR2[69] , 
        \Z\R_DATA_TEMPR3[69] , OR4_352_Y, \Z\R_DATA_TEMPR24[41] , 
        \Z\R_DATA_TEMPR25[41] , \Z\R_DATA_TEMPR26[41] , 
        \Z\R_DATA_TEMPR27[41] , OR4_153_Y, OR4_329_Y, OR4_400_Y, 
        OR4_470_Y, \Z\R_DATA_TEMPR28[53] , \Z\R_DATA_TEMPR29[53] , 
        \Z\R_DATA_TEMPR30[53] , \Z\R_DATA_TEMPR31[53] , OR4_456_Y, 
        \Z\R_DATA_TEMPR0[55] , \Z\R_DATA_TEMPR1[55] , 
        \Z\R_DATA_TEMPR2[55] , \Z\R_DATA_TEMPR3[55] , OR4_125_Y, 
        OR4_38_Y, OR4_425_Y, OR4_531_Y, OR4_636_Y, OR4_204_Y, 
        OR4_612_Y, OR4_646_Y, OR4_284_Y, \Z\R_DATA_TEMPR28[47] , 
        \Z\R_DATA_TEMPR29[47] , \Z\R_DATA_TEMPR30[47] , 
        \Z\R_DATA_TEMPR31[47] , \Z\R_DATA_TEMPR24[38] , 
        \Z\R_DATA_TEMPR25[38] , \Z\R_DATA_TEMPR26[38] , 
        \Z\R_DATA_TEMPR27[38] , \Z\R_DATA_TEMPR28[3] , 
        \Z\R_DATA_TEMPR29[3] , \Z\R_DATA_TEMPR30[3] , 
        \Z\R_DATA_TEMPR31[3] , \Z\R_DATA_TEMPR1[20] , 
        \Z\R_DATA_TEMPR1[21] , \Z\R_DATA_TEMPR1[23] , 
        \Z\R_DATA_TEMPR1[24] , \Z\R_DATA_TEMPR1[25] , 
        \Z\R_DATA_TEMPR1[27] , \Z\R_DATA_TEMPR1[28] , 
        \Z\R_DATA_TEMPR1[29] , \Z\R_DATA_TEMPR1[30] , 
        \Z\R_DATA_TEMPR1[31] , \Z\R_DATA_TEMPR1[35] , 
        \Z\R_DATA_TEMPR1[36] , \Z\R_DATA_TEMPR1[38] , 
        \Z\R_DATA_TEMPR1[39] , \Z\R_DATA_TEMPR1[1] , 
        \Z\R_DATA_TEMPR1[2] , \Z\R_DATA_TEMPR1[3] , 
        \Z\R_DATA_TEMPR1[4] , \Z\R_DATA_TEMPR1[6] , 
        \Z\R_DATA_TEMPR1[7] , \Z\R_DATA_TEMPR1[8] , 
        \Z\R_DATA_TEMPR1[9] , \Z\R_DATA_TEMPR1[11] , 
        \Z\R_DATA_TEMPR1[12] , \Z\R_DATA_TEMPR1[13] , 
        \Z\R_DATA_TEMPR1[14] , \Z\R_DATA_TEMPR1[15] , 
        \Z\R_DATA_TEMPR1[16] , \Z\R_DATA_TEMPR1[17] , 
        \Z\R_DATA_TEMPR1[18] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0_DB_DETECT, 
        \Z\ACCESS_BUSY[1][0] , OR4_588_Y, OR4_465_Y, OR4_396_Y, 
        \Z\R_DATA_TEMPR12[38] , \Z\R_DATA_TEMPR13[38] , 
        \Z\R_DATA_TEMPR14[38] , \Z\R_DATA_TEMPR15[38] , OR4_301_Y, 
        \Z\R_DATA_TEMPR24[20] , \Z\R_DATA_TEMPR25[20] , 
        \Z\R_DATA_TEMPR26[20] , \Z\R_DATA_TEMPR27[20] , OR4_95_Y, 
        OR4_385_Y, OR4_5_Y, OR4_55_Y, \Z\R_DATA_TEMPR12[57] , 
        \Z\R_DATA_TEMPR13[57] , \Z\R_DATA_TEMPR15[57] , OR4_558_Y, 
        OR4_188_Y, OR4_687_Y, OR4_1_Y, OR4_494_Y, 
        \Z\R_DATA_TEMPR28[35] , \Z\R_DATA_TEMPR29[35] , 
        \Z\R_DATA_TEMPR30[35] , \Z\R_DATA_TEMPR31[35] , OR2_11_Y, 
        \Z\R_DATA_TEMPR21[50] , \Z\R_DATA_TEMPR8[48] , 
        \Z\R_DATA_TEMPR9[48] , \Z\R_DATA_TEMPR10[48] , 
        \Z\R_DATA_TEMPR11[48] , OR4_504_Y, OR4_121_Y, OR4_73_Y, 
        \Z\R_DATA_TEMPR4[15] , \Z\R_DATA_TEMPR6[15] , 
        \Z\R_DATA_TEMPR7[15] , OR4_142_Y, \Z\R_DATA_TEMPR24[31] , 
        \Z\R_DATA_TEMPR25[31] , \Z\R_DATA_TEMPR26[31] , 
        \Z\R_DATA_TEMPR27[31] , OR4_154_Y, OR4_501_Y, OR4_29_Y, 
        OR2_71_Y, \Z\R_DATA_TEMPR21[27] , OR4_618_Y, 
        \Z\R_DATA_TEMPR24[62] , \Z\R_DATA_TEMPR25[62] , 
        \Z\R_DATA_TEMPR26[62] , \Z\R_DATA_TEMPR27[62] , OR2_54_Y, 
        \Z\R_DATA_TEMPR21[59] , \Z\R_DATA_TEMPR0[14] , 
        \Z\R_DATA_TEMPR2[14] , \Z\R_DATA_TEMPR3[14] , OR4_495_Y, 
        OR4_626_Y, OR4_486_Y, OR4_108_Y, OR4_556_Y, OR4_78_Y, 
        OR4_225_Y, OR4_86_Y, OR4_463_Y, OR4_233_Y, OR4_350_Y, 
        OR4_388_Y, OR4_502_Y, OR4_209_Y, \Z\R_DATA_TEMPR22[12] , 
        \Z\R_DATA_TEMPR28[20] , \Z\R_DATA_TEMPR28[21] , 
        \Z\R_DATA_TEMPR28[22] , \Z\R_DATA_TEMPR28[25] , 
        \Z\R_DATA_TEMPR28[27] , \Z\R_DATA_TEMPR28[29] , 
        \Z\R_DATA_TEMPR28[30] , \Z\R_DATA_TEMPR28[31] , 
        \Z\R_DATA_TEMPR28[32] , \Z\R_DATA_TEMPR28[33] , 
        \Z\R_DATA_TEMPR28[36] , \Z\R_DATA_TEMPR28[37] , 
        \Z\R_DATA_TEMPR28[38] , \Z\R_DATA_TEMPR28[39] , 
        \Z\R_DATA_TEMPR28[1] , \Z\R_DATA_TEMPR28[2] , 
        \Z\R_DATA_TEMPR28[4] , \Z\R_DATA_TEMPR28[5] , 
        \Z\R_DATA_TEMPR28[6] , \Z\R_DATA_TEMPR28[7] , 
        \Z\R_DATA_TEMPR28[8] , \Z\R_DATA_TEMPR28[10] , 
        \Z\R_DATA_TEMPR28[11] , \Z\R_DATA_TEMPR28[12] , 
        \Z\R_DATA_TEMPR28[13] , \Z\R_DATA_TEMPR28[14] , 
        \Z\R_DATA_TEMPR28[15] , \Z\R_DATA_TEMPR28[16] , 
        \Z\R_DATA_TEMPR28[17] , \Z\R_DATA_TEMPR28[18] , 
        \Z\R_DATA_TEMPR28[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0_DB_DETECT, 
        \Z\ACCESS_BUSY[28][0] , OR4_460_Y, \Z\R_DATA_TEMPR12[63] , 
        \Z\R_DATA_TEMPR13[63] , \Z\R_DATA_TEMPR15[63] , 
        \Z\R_DATA_TEMPR24[60] , \Z\R_DATA_TEMPR24[61] , 
        \Z\R_DATA_TEMPR24[63] , \Z\R_DATA_TEMPR24[65] , 
        \Z\R_DATA_TEMPR24[66] , \Z\R_DATA_TEMPR24[67] , 
        \Z\R_DATA_TEMPR24[68] , \Z\R_DATA_TEMPR24[69] , 
        \Z\R_DATA_TEMPR24[70] , \Z\R_DATA_TEMPR24[71] , 
        \Z\R_DATA_TEMPR24[72] , \Z\R_DATA_TEMPR24[73] , 
        \Z\R_DATA_TEMPR24[74] , \Z\R_DATA_TEMPR24[75] , 
        \Z\R_DATA_TEMPR24[77] , \Z\R_DATA_TEMPR24[78] , 
        \Z\R_DATA_TEMPR24[79] , \Z\R_DATA_TEMPR24[40] , 
        \Z\R_DATA_TEMPR24[42] , \Z\R_DATA_TEMPR24[43] , 
        \Z\R_DATA_TEMPR24[44] , \Z\R_DATA_TEMPR24[47] , 
        \Z\R_DATA_TEMPR24[48] , \Z\R_DATA_TEMPR24[49] , 
        \Z\R_DATA_TEMPR24[50] , \Z\R_DATA_TEMPR24[51] , 
        \Z\R_DATA_TEMPR24[52] , \Z\R_DATA_TEMPR24[53] , 
        \Z\R_DATA_TEMPR24[54] , \Z\R_DATA_TEMPR24[55] , 
        \Z\R_DATA_TEMPR24[57] , \Z\R_DATA_TEMPR24[58] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C1_DB_DETECT, 
        \Z\ACCESS_BUSY[24][1] , OR4_271_Y, \Z\R_DATA_TEMPR4[45] , 
        \Z\R_DATA_TEMPR5[45] , \Z\R_DATA_TEMPR7[45] , OR4_6_Y, 
        OR4_182_Y, OR2_67_Y, \Z\R_DATA_TEMPR22[16] , 
        \Z\R_DATA_TEMPR21[20] , \Z\R_DATA_TEMPR21[21] , 
        \Z\R_DATA_TEMPR21[22] , \Z\R_DATA_TEMPR21[23] , 
        \Z\R_DATA_TEMPR21[24] , \Z\R_DATA_TEMPR21[25] , 
        \Z\R_DATA_TEMPR21[26] , \Z\R_DATA_TEMPR21[28] , 
        \Z\R_DATA_TEMPR21[29] , \Z\R_DATA_TEMPR21[31] , 
        \Z\R_DATA_TEMPR21[32] , \Z\R_DATA_TEMPR21[34] , 
        \Z\R_DATA_TEMPR21[35] , \Z\R_DATA_TEMPR21[36] , 
        \Z\R_DATA_TEMPR21[37] , \Z\R_DATA_TEMPR21[38] , 
        \Z\R_DATA_TEMPR21[39] , \Z\R_DATA_TEMPR21[0] , 
        \Z\R_DATA_TEMPR21[1] , \Z\R_DATA_TEMPR21[2] , 
        \Z\R_DATA_TEMPR21[3] , \Z\R_DATA_TEMPR21[4] , 
        \Z\R_DATA_TEMPR21[5] , \Z\R_DATA_TEMPR21[6] , 
        \Z\R_DATA_TEMPR21[7] , \Z\R_DATA_TEMPR21[8] , 
        \Z\R_DATA_TEMPR21[10] , \Z\R_DATA_TEMPR21[11] , 
        \Z\R_DATA_TEMPR21[16] , \Z\R_DATA_TEMPR21[17] , 
        \Z\R_DATA_TEMPR21[18] , \Z\R_DATA_TEMPR21[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0_DB_DETECT, 
        \Z\ACCESS_BUSY[21][0] , OR4_81_Y, OR4_578_Y, OR4_299_Y, 
        OR4_660_Y, OR4_402_Y, OR4_39_Y, OR4_348_Y, OR4_361_Y, 
        \Z\R_DATA_TEMPR29[18] , \Z\R_DATA_TEMPR30[18] , 
        \Z\R_DATA_TEMPR31[18] , OR4_201_Y, \Z\R_DATA_TEMPR4[43] , 
        \Z\R_DATA_TEMPR5[43] , \Z\R_DATA_TEMPR7[43] , OR4_213_Y, 
        \Z\R_DATA_TEMPR25[73] , \Z\R_DATA_TEMPR26[73] , 
        \Z\R_DATA_TEMPR27[73] , OR4_632_Y, \Z\R_DATA_TEMPR25[50] , 
        \Z\R_DATA_TEMPR26[50] , \Z\R_DATA_TEMPR27[50] , OR4_143_Y, 
        \Z\R_DATA_TEMPR12[8] , \Z\R_DATA_TEMPR13[8] , 
        \Z\R_DATA_TEMPR14[8] , \Z\R_DATA_TEMPR15[8] , 
        \Z\R_DATA_TEMPR29[20] , \Z\R_DATA_TEMPR29[21] , 
        \Z\R_DATA_TEMPR29[22] , \Z\R_DATA_TEMPR29[25] , 
        \Z\R_DATA_TEMPR29[27] , \Z\R_DATA_TEMPR29[29] , 
        \Z\R_DATA_TEMPR29[30] , \Z\R_DATA_TEMPR29[31] , 
        \Z\R_DATA_TEMPR29[32] , \Z\R_DATA_TEMPR29[33] , 
        \Z\R_DATA_TEMPR29[36] , \Z\R_DATA_TEMPR29[37] , 
        \Z\R_DATA_TEMPR29[38] , \Z\R_DATA_TEMPR29[39] , 
        \Z\R_DATA_TEMPR29[1] , \Z\R_DATA_TEMPR29[2] , 
        \Z\R_DATA_TEMPR29[4] , \Z\R_DATA_TEMPR29[5] , 
        \Z\R_DATA_TEMPR29[6] , \Z\R_DATA_TEMPR29[7] , 
        \Z\R_DATA_TEMPR29[8] , \Z\R_DATA_TEMPR29[10] , 
        \Z\R_DATA_TEMPR29[11] , \Z\R_DATA_TEMPR29[12] , 
        \Z\R_DATA_TEMPR29[13] , \Z\R_DATA_TEMPR29[14] , 
        \Z\R_DATA_TEMPR29[15] , \Z\R_DATA_TEMPR29[16] , 
        \Z\R_DATA_TEMPR29[17] , \Z\R_DATA_TEMPR29[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0_DB_DETECT, 
        \Z\ACCESS_BUSY[29][0] , \Z\R_DATA_TEMPR21[75] , OR4_22_Y, 
        \Z\R_DATA_TEMPR8[41] , \Z\R_DATA_TEMPR9[41] , 
        \Z\R_DATA_TEMPR10[41] , \Z\R_DATA_TEMPR11[41] , OR4_638_Y, 
        \Z\R_DATA_TEMPR0[38] , \Z\R_DATA_TEMPR2[38] , 
        \Z\R_DATA_TEMPR3[38] , OR2_21_Y, OR4_684_Y, 
        \Z\R_DATA_TEMPR0[16] , \Z\R_DATA_TEMPR2[16] , 
        \Z\R_DATA_TEMPR3[16] , OR4_230_Y, OR4_193_Y, OR4_210_Y, 
        OR4_697_Y, OR4_223_Y, OR4_614_Y, OR4_167_Y, OR4_512_Y, 
        OR4_564_Y, OR4_190_Y, OR2_1_Y, \Z\R_DATA_TEMPR22[78] , 
        \Z\R_DATA_TEMPR23[78] , OR4_362_Y, OR4_441_Y, OR4_275_Y, 
        OR4_542_Y, OR4_403_Y, OR4_10_Y, OR4_454_Y, 
        \Z\R_DATA_TEMPR0[4] , \Z\R_DATA_TEMPR2[4] , 
        \Z\R_DATA_TEMPR3[4] , OR4_286_Y, OR2_7_Y, 
        \Z\R_DATA_TEMPR22[69] , \Z\R_DATA_TEMPR23[69] , 
        \Z\R_DATA_TEMPR12[20] , \Z\R_DATA_TEMPR12[21] , 
        \Z\R_DATA_TEMPR12[22] , \Z\R_DATA_TEMPR12[23] , 
        \Z\R_DATA_TEMPR12[24] , \Z\R_DATA_TEMPR12[28] , 
        \Z\R_DATA_TEMPR12[29] , \Z\R_DATA_TEMPR12[30] , 
        \Z\R_DATA_TEMPR12[31] , \Z\R_DATA_TEMPR12[32] , 
        \Z\R_DATA_TEMPR12[33] , \Z\R_DATA_TEMPR12[35] , 
        \Z\R_DATA_TEMPR12[36] , \Z\R_DATA_TEMPR12[39] , 
        \Z\R_DATA_TEMPR12[0] , \Z\R_DATA_TEMPR12[1] , 
        \Z\R_DATA_TEMPR12[2] , \Z\R_DATA_TEMPR12[3] , 
        \Z\R_DATA_TEMPR12[4] , \Z\R_DATA_TEMPR12[5] , 
        \Z\R_DATA_TEMPR12[6] , \Z\R_DATA_TEMPR12[7] , 
        \Z\R_DATA_TEMPR12[9] , \Z\R_DATA_TEMPR12[10] , 
        \Z\R_DATA_TEMPR12[11] , \Z\R_DATA_TEMPR12[13] , 
        \Z\R_DATA_TEMPR12[14] , \Z\R_DATA_TEMPR12[15] , 
        \Z\R_DATA_TEMPR12[16] , \Z\R_DATA_TEMPR12[17] , 
        \Z\R_DATA_TEMPR12[18] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0_DB_DETECT, 
        \Z\ACCESS_BUSY[12][0] , OR4_643_Y, \Z\R_DATA_TEMPR4[51] , 
        \Z\R_DATA_TEMPR5[51] , \Z\R_DATA_TEMPR7[51] , OR4_689_Y, 
        OR4_467_Y, OR4_212_Y, OR4_244_Y, \Z\R_DATA_TEMPR3[20] , 
        \Z\R_DATA_TEMPR3[21] , \Z\R_DATA_TEMPR3[23] , 
        \Z\R_DATA_TEMPR3[24] , \Z\R_DATA_TEMPR3[25] , 
        \Z\R_DATA_TEMPR3[27] , \Z\R_DATA_TEMPR3[28] , 
        \Z\R_DATA_TEMPR3[29] , \Z\R_DATA_TEMPR3[30] , 
        \Z\R_DATA_TEMPR3[31] , \Z\R_DATA_TEMPR3[35] , 
        \Z\R_DATA_TEMPR3[36] , \Z\R_DATA_TEMPR3[39] , 
        \Z\R_DATA_TEMPR3[1] , \Z\R_DATA_TEMPR3[2] , 
        \Z\R_DATA_TEMPR3[3] , \Z\R_DATA_TEMPR3[6] , 
        \Z\R_DATA_TEMPR3[7] , \Z\R_DATA_TEMPR3[8] , 
        \Z\R_DATA_TEMPR3[9] , \Z\R_DATA_TEMPR3[11] , 
        \Z\R_DATA_TEMPR3[12] , \Z\R_DATA_TEMPR3[13] , 
        \Z\R_DATA_TEMPR3[15] , \Z\R_DATA_TEMPR3[17] , 
        \Z\R_DATA_TEMPR3[18] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0_DB_DETECT, 
        \Z\ACCESS_BUSY[3][0] , OR4_506_Y, OR4_513_Y, OR4_109_Y, 
        OR4_378_Y, OR4_341_Y, OR4_120_Y, OR4_390_Y, 
        \Z\R_DATA_TEMPR22[66] , \Z\R_DATA_TEMPR23[66] , 
        \Z\R_DATA_TEMPR8[47] , \Z\R_DATA_TEMPR9[47] , 
        \Z\R_DATA_TEMPR10[47] , \Z\R_DATA_TEMPR11[47] , 
        \Z\R_DATA_TEMPR27[60] , \Z\R_DATA_TEMPR27[61] , 
        \Z\R_DATA_TEMPR27[63] , \Z\R_DATA_TEMPR27[65] , 
        \Z\R_DATA_TEMPR27[66] , \Z\R_DATA_TEMPR27[67] , 
        \Z\R_DATA_TEMPR27[68] , \Z\R_DATA_TEMPR27[69] , 
        \Z\R_DATA_TEMPR27[70] , \Z\R_DATA_TEMPR27[71] , 
        \Z\R_DATA_TEMPR27[72] , \Z\R_DATA_TEMPR27[74] , 
        \Z\R_DATA_TEMPR27[75] , \Z\R_DATA_TEMPR27[77] , 
        \Z\R_DATA_TEMPR27[78] , \Z\R_DATA_TEMPR27[79] , 
        \Z\R_DATA_TEMPR27[40] , \Z\R_DATA_TEMPR27[42] , 
        \Z\R_DATA_TEMPR27[43] , \Z\R_DATA_TEMPR27[44] , 
        \Z\R_DATA_TEMPR27[47] , \Z\R_DATA_TEMPR27[48] , 
        \Z\R_DATA_TEMPR27[49] , \Z\R_DATA_TEMPR27[51] , 
        \Z\R_DATA_TEMPR27[52] , \Z\R_DATA_TEMPR27[53] , 
        \Z\R_DATA_TEMPR27[54] , \Z\R_DATA_TEMPR27[55] , 
        \Z\R_DATA_TEMPR27[57] , \Z\R_DATA_TEMPR27[58] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C1_DB_DETECT, 
        \Z\ACCESS_BUSY[27][1] , OR4_587_Y, \Z\R_DATA_TEMPR19[48] , 
        OR4_280_Y, OR4_407_Y, OR4_330_Y, OR4_129_Y, OR4_173_Y, 
        \Z\R_DATA_TEMPR30[17] , \Z\R_DATA_TEMPR31[17] , OR2_23_Y, 
        \Z\R_DATA_TEMPR21[77] , OR4_261_Y, \Z\R_DATA_TEMPR25[51] , 
        \Z\R_DATA_TEMPR26[51] , \Z\R_DATA_TEMPR4[12] , 
        \Z\R_DATA_TEMPR6[12] , \Z\R_DATA_TEMPR7[12] , OR4_229_Y, 
        \Z\R_DATA_TEMPR0[71] , \Z\R_DATA_TEMPR1[71] , 
        \Z\R_DATA_TEMPR2[71] , \Z\R_DATA_TEMPR3[71] , OR4_593_Y, 
        OR4_34_Y, OR4_76_Y, OR4_67_Y, OR4_701_Y, 
        \Z\R_DATA_TEMPR28[40] , \Z\R_DATA_TEMPR29[40] , 
        \Z\R_DATA_TEMPR30[40] , \Z\R_DATA_TEMPR31[40] , 
        \Z\R_DATA_TEMPR0[20] , \Z\R_DATA_TEMPR0[21] , 
        \Z\R_DATA_TEMPR0[23] , \Z\R_DATA_TEMPR0[24] , 
        \Z\R_DATA_TEMPR0[25] , \Z\R_DATA_TEMPR0[27] , 
        \Z\R_DATA_TEMPR0[28] , \Z\R_DATA_TEMPR0[29] , 
        \Z\R_DATA_TEMPR0[30] , \Z\R_DATA_TEMPR0[31] , 
        \Z\R_DATA_TEMPR0[35] , \Z\R_DATA_TEMPR0[36] , 
        \Z\R_DATA_TEMPR0[39] , \Z\R_DATA_TEMPR0[1] , 
        \Z\R_DATA_TEMPR0[2] , \Z\R_DATA_TEMPR0[3] , 
        \Z\R_DATA_TEMPR0[6] , \Z\R_DATA_TEMPR0[7] , 
        \Z\R_DATA_TEMPR0[8] , \Z\R_DATA_TEMPR0[9] , 
        \Z\R_DATA_TEMPR0[11] , \Z\R_DATA_TEMPR0[12] , 
        \Z\R_DATA_TEMPR0[13] , \Z\R_DATA_TEMPR0[15] , 
        \Z\R_DATA_TEMPR0[17] , \Z\R_DATA_TEMPR0[18] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0_DB_DETECT, 
        \Z\ACCESS_BUSY[0][0] , OR4_138_Y, OR2_12_Y, 
        \Z\R_DATA_TEMPR22[10] , \Z\R_DATA_TEMPR8[70] , 
        \Z\R_DATA_TEMPR9[70] , \Z\R_DATA_TEMPR10[70] , 
        \Z\R_DATA_TEMPR11[70] , OR4_18_Y, \Z\R_DATA_TEMPR30[22] , 
        \Z\R_DATA_TEMPR31[22] , OR4_242_Y, OR4_417_Y, OR4_382_Y, 
        \Z\R_DATA_TEMPR4[10] , \Z\R_DATA_TEMPR6[10] , 
        \Z\R_DATA_TEMPR7[10] , OR4_122_Y, OR4_259_Y, OR4_2_Y, 
        OR4_691_Y, OR4_706_Y, OR4_481_Y, \Z\R_DATA_TEMPR26[60] , 
        \Z\R_DATA_TEMPR26[61] , \Z\R_DATA_TEMPR26[63] , 
        \Z\R_DATA_TEMPR26[65] , \Z\R_DATA_TEMPR26[66] , 
        \Z\R_DATA_TEMPR26[67] , \Z\R_DATA_TEMPR26[68] , 
        \Z\R_DATA_TEMPR26[69] , \Z\R_DATA_TEMPR26[70] , 
        \Z\R_DATA_TEMPR26[71] , \Z\R_DATA_TEMPR26[72] , 
        \Z\R_DATA_TEMPR26[74] , \Z\R_DATA_TEMPR26[75] , 
        \Z\R_DATA_TEMPR26[77] , \Z\R_DATA_TEMPR26[78] , 
        \Z\R_DATA_TEMPR26[79] , \Z\R_DATA_TEMPR26[40] , 
        \Z\R_DATA_TEMPR26[42] , \Z\R_DATA_TEMPR26[43] , 
        \Z\R_DATA_TEMPR26[44] , \Z\R_DATA_TEMPR26[47] , 
        \Z\R_DATA_TEMPR26[48] , \Z\R_DATA_TEMPR26[49] , 
        \Z\R_DATA_TEMPR26[52] , \Z\R_DATA_TEMPR26[53] , 
        \Z\R_DATA_TEMPR26[54] , \Z\R_DATA_TEMPR26[55] , 
        \Z\R_DATA_TEMPR26[57] , \Z\R_DATA_TEMPR26[58] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C1_DB_DETECT, 
        \Z\ACCESS_BUSY[26][1] , OR4_719_Y, \Z\R_DATA_TEMPR8[49] , 
        \Z\R_DATA_TEMPR9[49] , \Z\R_DATA_TEMPR10[49] , 
        \Z\R_DATA_TEMPR11[49] , OR4_340_Y, \Z\R_DATA_TEMPR16[36] , 
        \Z\R_DATA_TEMPR17[36] , OR2_52_Y, OR4_107_Y, OR4_457_Y, 
        OR4_601_Y, \Z\R_DATA_TEMPR8[72] , \Z\R_DATA_TEMPR9[72] , 
        \Z\R_DATA_TEMPR10[72] , \Z\R_DATA_TEMPR11[72] , OR4_455_Y, 
        \Z\R_DATA_TEMPR12[71] , \Z\R_DATA_TEMPR13[71] , 
        \Z\R_DATA_TEMPR15[71] , \Z\R_DATA_TEMPR25[71] , 
        \Z\R_DATA_TEMPR28[60] , \Z\R_DATA_TEMPR29[60] , 
        \Z\R_DATA_TEMPR30[60] , \Z\R_DATA_TEMPR31[60] , OR4_604_Y, 
        OR4_65_Y, OR2_36_Y, \Z\R_DATA_TEMPR22[34] , OR4_77_Y, 
        \Z\R_DATA_TEMPR8[35] , OR4_375_Y, \Z\R_DATA_TEMPR22[9] , 
        OR4_276_Y, \Z\R_DATA_TEMPR4[54] , \Z\R_DATA_TEMPR5[54] , 
        \Z\R_DATA_TEMPR7[54] , \Z\R_DATA_TEMPR30[39] , 
        \Z\R_DATA_TEMPR31[39] , \Z\R_DATA_TEMPR4[58] , 
        \Z\R_DATA_TEMPR5[58] , \Z\R_DATA_TEMPR7[58] , 
        \Z\R_DATA_TEMPR25[55] , OR4_533_Y, \Z\R_DATA_TEMPR8[7] , 
        OR4_206_Y, OR4_57_Y, OR2_24_Y, \Z\R_DATA_TEMPR22[23] , 
        \Z\R_DATA_TEMPR14[20] , \Z\R_DATA_TEMPR14[21] , 
        \Z\R_DATA_TEMPR14[22] , \Z\R_DATA_TEMPR14[23] , 
        \Z\R_DATA_TEMPR14[24] , \Z\R_DATA_TEMPR14[28] , 
        \Z\R_DATA_TEMPR14[29] , \Z\R_DATA_TEMPR14[30] , 
        \Z\R_DATA_TEMPR14[31] , \Z\R_DATA_TEMPR14[32] , 
        \Z\R_DATA_TEMPR14[33] , \Z\R_DATA_TEMPR14[35] , 
        \Z\R_DATA_TEMPR14[36] , \Z\R_DATA_TEMPR14[39] , 
        \Z\R_DATA_TEMPR14[0] , \Z\R_DATA_TEMPR14[1] , 
        \Z\R_DATA_TEMPR14[2] , \Z\R_DATA_TEMPR14[3] , 
        \Z\R_DATA_TEMPR14[4] , \Z\R_DATA_TEMPR14[5] , 
        \Z\R_DATA_TEMPR14[6] , \Z\R_DATA_TEMPR14[7] , 
        \Z\R_DATA_TEMPR14[9] , \Z\R_DATA_TEMPR14[10] , 
        \Z\R_DATA_TEMPR14[11] , \Z\R_DATA_TEMPR14[13] , 
        \Z\R_DATA_TEMPR14[14] , \Z\R_DATA_TEMPR14[15] , 
        \Z\R_DATA_TEMPR14[16] , \Z\R_DATA_TEMPR14[17] , 
        \Z\R_DATA_TEMPR14[18] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0_DB_DETECT, 
        \Z\ACCESS_BUSY[14][0] , OR4_679_Y, \Z\R_DATA_TEMPR2[13] , 
        OR4_123_Y, \Z\R_DATA_TEMPR2[25] , \Z\R_DATA_TEMPR28[61] , 
        \Z\R_DATA_TEMPR28[62] , \Z\R_DATA_TEMPR28[63] , 
        \Z\R_DATA_TEMPR28[66] , \Z\R_DATA_TEMPR28[67] , 
        \Z\R_DATA_TEMPR28[68] , \Z\R_DATA_TEMPR28[69] , 
        \Z\R_DATA_TEMPR28[71] , \Z\R_DATA_TEMPR28[72] , 
        \Z\R_DATA_TEMPR28[73] , \Z\R_DATA_TEMPR28[74] , 
        \Z\R_DATA_TEMPR28[75] , \Z\R_DATA_TEMPR28[76] , 
        \Z\R_DATA_TEMPR28[77] , \Z\R_DATA_TEMPR28[79] , 
        \Z\R_DATA_TEMPR28[41] , \Z\R_DATA_TEMPR28[42] , 
        \Z\R_DATA_TEMPR28[43] , \Z\R_DATA_TEMPR28[44] , 
        \Z\R_DATA_TEMPR28[45] , \Z\R_DATA_TEMPR28[48] , 
        \Z\R_DATA_TEMPR28[49] , \Z\R_DATA_TEMPR28[50] , 
        \Z\R_DATA_TEMPR28[51] , \Z\R_DATA_TEMPR28[52] , 
        \Z\R_DATA_TEMPR28[54] , \Z\R_DATA_TEMPR28[57] , 
        \Z\R_DATA_TEMPR28[58] , \Z\R_DATA_TEMPR28[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C1_DB_DETECT, 
        \Z\ACCESS_BUSY[28][1] , \Z\R_DATA_TEMPR12[48] , 
        \Z\R_DATA_TEMPR13[48] , \Z\R_DATA_TEMPR15[48] , OR4_319_Y, 
        \Z\R_DATA_TEMPR16[29] , \Z\R_DATA_TEMPR17[29] , 
        \Z\R_DATA_TEMPR12[56] , \Z\R_DATA_TEMPR13[56] , 
        \Z\R_DATA_TEMPR15[56] , OR4_541_Y, \Z\R_DATA_TEMPR4[13] , 
        \Z\R_DATA_TEMPR6[13] , \Z\R_DATA_TEMPR7[13] , OR4_577_Y, 
        \Z\R_DATA_TEMPR29[43] , \Z\R_DATA_TEMPR30[43] , 
        \Z\R_DATA_TEMPR31[43] , \Z\R_DATA_TEMPR12[44] , 
        \Z\R_DATA_TEMPR13[44] , \Z\R_DATA_TEMPR15[44] , 
        \Z\R_DATA_TEMPR21[46] , \Z\R_DATA_TEMPR4[73] , 
        \Z\R_DATA_TEMPR5[73] , \Z\R_DATA_TEMPR7[73] , OR4_189_Y, 
        OR4_652_Y, OR4_200_Y, \Z\R_DATA_TEMPR2[21] , OR4_586_Y, 
        \Z\R_DATA_TEMPR8[61] , \Z\R_DATA_TEMPR9[61] , 
        \Z\R_DATA_TEMPR10[61] , \Z\R_DATA_TEMPR11[61] , OR4_623_Y, 
        \Z\R_DATA_TEMPR0[41] , \Z\R_DATA_TEMPR1[41] , 
        \Z\R_DATA_TEMPR2[41] , \Z\R_DATA_TEMPR3[41] , 
        \Z\R_DATA_TEMPR13[67] , \Z\R_DATA_TEMPR13[69] , 
        \Z\R_DATA_TEMPR13[70] , \Z\R_DATA_TEMPR13[72] , 
        \Z\R_DATA_TEMPR13[73] , \Z\R_DATA_TEMPR13[74] , 
        \Z\R_DATA_TEMPR13[75] , \Z\R_DATA_TEMPR13[76] , 
        \Z\R_DATA_TEMPR13[77] , \Z\R_DATA_TEMPR13[40] , 
        \Z\R_DATA_TEMPR13[41] , \Z\R_DATA_TEMPR13[43] , 
        \Z\R_DATA_TEMPR13[45] , \Z\R_DATA_TEMPR13[46] , 
        \Z\R_DATA_TEMPR13[47] , \Z\R_DATA_TEMPR13[50] , 
        \Z\R_DATA_TEMPR13[51] , \Z\R_DATA_TEMPR13[53] , 
        \Z\R_DATA_TEMPR13[54] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C1_DB_DETECT, 
        \Z\ACCESS_BUSY[13][1] , OR4_150_Y, \Z\R_DATA_TEMPR22[71] , 
        \Z\R_DATA_TEMPR23[71] , \Z\R_DATA_TEMPR4[56] , 
        \Z\R_DATA_TEMPR5[56] , \Z\R_DATA_TEMPR7[56] , OR4_525_Y, 
        \Z\R_DATA_TEMPR8[0] , OR4_84_Y, OR4_430_Y, OR4_32_Y, OR4_372_Y, 
        \Z\R_DATA_TEMPR25[72] , \Z\R_DATA_TEMPR4[60] , 
        \Z\R_DATA_TEMPR4[61] , \Z\R_DATA_TEMPR4[62] , 
        \Z\R_DATA_TEMPR4[63] , \Z\R_DATA_TEMPR4[65] , 
        \Z\R_DATA_TEMPR4[66] , \Z\R_DATA_TEMPR4[67] , 
        \Z\R_DATA_TEMPR4[68] , \Z\R_DATA_TEMPR4[69] , 
        \Z\R_DATA_TEMPR4[78] , \Z\R_DATA_TEMPR4[79] , 
        \Z\R_DATA_TEMPR4[40] , \Z\R_DATA_TEMPR4[41] , 
        \Z\R_DATA_TEMPR4[44] , \Z\R_DATA_TEMPR4[46] , 
        \Z\R_DATA_TEMPR4[49] , \Z\R_DATA_TEMPR4[50] , 
        \Z\R_DATA_TEMPR4[52] , \Z\R_DATA_TEMPR4[55] , 
        \Z\R_DATA_TEMPR4[57] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C1_DB_DETECT, 
        \Z\ACCESS_BUSY[4][1] , OR4_394_Y, OR2_63_Y, 
        \Z\R_DATA_TEMPR22[61] , \Z\R_DATA_TEMPR23[61] , OR4_339_Y, 
        \Z\R_DATA_TEMPR24[22] , \Z\R_DATA_TEMPR25[22] , 
        \Z\R_DATA_TEMPR26[22] , \Z\R_DATA_TEMPR27[22] , OR4_410_Y, 
        \Z\R_DATA_TEMPR5[49] , \Z\R_DATA_TEMPR7[49] , 
        \Z\R_DATA_TEMPR30[10] , \Z\R_DATA_TEMPR31[10] , OR4_25_Y, 
        \Z\R_DATA_TEMPR29[51] , \Z\R_DATA_TEMPR30[51] , 
        \Z\R_DATA_TEMPR31[51] , \Z\R_DATA_TEMPR25[40] , 
        \Z\R_DATA_TEMPR8[60] , \Z\R_DATA_TEMPR8[62] , 
        \Z\R_DATA_TEMPR8[63] , \Z\R_DATA_TEMPR8[64] , 
        \Z\R_DATA_TEMPR8[65] , \Z\R_DATA_TEMPR8[66] , 
        \Z\R_DATA_TEMPR8[67] , \Z\R_DATA_TEMPR8[68] , 
        \Z\R_DATA_TEMPR8[69] , \Z\R_DATA_TEMPR8[73] , 
        \Z\R_DATA_TEMPR8[74] , \Z\R_DATA_TEMPR8[76] , 
        \Z\R_DATA_TEMPR8[40] , \Z\R_DATA_TEMPR8[42] , 
        \Z\R_DATA_TEMPR8[43] , \Z\R_DATA_TEMPR8[44] , 
        \Z\R_DATA_TEMPR8[46] , \Z\R_DATA_TEMPR8[51] , 
        \Z\R_DATA_TEMPR8[52] , \Z\R_DATA_TEMPR8[53] , 
        \Z\R_DATA_TEMPR8[55] , \Z\R_DATA_TEMPR8[57] , 
        \Z\R_DATA_TEMPR8[58] , \Z\R_DATA_TEMPR8[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C1_DB_DETECT, 
        \Z\ACCESS_BUSY[8][1] , OR4_266_Y, OR4_113_Y, 
        \Z\R_DATA_TEMPR22[13] , OR4_302_Y, \Z\R_DATA_TEMPR24[36] , 
        \Z\R_DATA_TEMPR25[36] , \Z\R_DATA_TEMPR26[36] , 
        \Z\R_DATA_TEMPR27[36] , OR4_248_Y, \Z\R_DATA_TEMPR25[78] , 
        OR4_311_Y, \Z\R_DATA_TEMPR13[30] , \Z\R_DATA_TEMPR15[30] , 
        OR4_184_Y, \Z\R_DATA_TEMPR0[63] , \Z\R_DATA_TEMPR1[63] , 
        \Z\R_DATA_TEMPR2[63] , \Z\R_DATA_TEMPR3[63] , OR4_476_Y, 
        OR4_165_Y, OR2_64_Y, \Z\R_DATA_TEMPR22[72] , 
        \Z\R_DATA_TEMPR23[72] , OR4_641_Y, \Z\R_DATA_TEMPR25[48] , 
        OR4_669_Y, OR4_308_Y, OR4_307_Y, OR4_423_Y, OR4_443_Y, 
        \Z\R_DATA_TEMPR13[7] , \Z\R_DATA_TEMPR15[7] , OR4_406_Y, 
        \Z\R_DATA_TEMPR19[50] , \Z\R_DATA_TEMPR24[32] , 
        \Z\R_DATA_TEMPR25[32] , \Z\R_DATA_TEMPR26[32] , 
        \Z\R_DATA_TEMPR27[32] , OR4_260_Y, \Z\R_DATA_TEMPR13[13] , 
        \Z\R_DATA_TEMPR15[13] , \Z\R_DATA_TEMPR29[44] , 
        \Z\R_DATA_TEMPR30[44] , \Z\R_DATA_TEMPR31[44] , 
        \Z\R_DATA_TEMPR16[23] , \Z\R_DATA_TEMPR17[23] , OR4_693_Y, 
        \Z\R_DATA_TEMPR8[33] , \Z\R_DATA_TEMPR25[60] , 
        \Z\R_DATA_TEMPR12[53] , \Z\R_DATA_TEMPR15[53] , OR4_50_Y, 
        \Z\R_DATA_TEMPR4[35] , \Z\R_DATA_TEMPR6[35] , 
        \Z\R_DATA_TEMPR7[35] , \Z\R_DATA_TEMPR8[12] , 
        \Z\R_DATA_TEMPR0[56] , \Z\R_DATA_TEMPR1[56] , 
        \Z\R_DATA_TEMPR2[56] , \Z\R_DATA_TEMPR3[56] , OR4_595_Y, 
        \Z\R_DATA_TEMPR29[79] , \Z\R_DATA_TEMPR30[79] , 
        \Z\R_DATA_TEMPR31[79] , OR4_428_Y, OR4_60_Y, OR4_380_Y, 
        \Z\R_DATA_TEMPR7[20] , \Z\R_DATA_TEMPR7[21] , 
        \Z\R_DATA_TEMPR7[22] , \Z\R_DATA_TEMPR7[23] , 
        \Z\R_DATA_TEMPR7[26] , \Z\R_DATA_TEMPR7[28] , 
        \Z\R_DATA_TEMPR7[29] , \Z\R_DATA_TEMPR7[30] , 
        \Z\R_DATA_TEMPR7[31] , \Z\R_DATA_TEMPR7[37] , 
        \Z\R_DATA_TEMPR7[38] , \Z\R_DATA_TEMPR7[0] , 
        \Z\R_DATA_TEMPR7[1] , \Z\R_DATA_TEMPR7[2] , 
        \Z\R_DATA_TEMPR7[3] , \Z\R_DATA_TEMPR7[4] , 
        \Z\R_DATA_TEMPR7[5] , \Z\R_DATA_TEMPR7[6] , 
        \Z\R_DATA_TEMPR7[8] , \Z\R_DATA_TEMPR7[9] , 
        \Z\R_DATA_TEMPR7[14] , \Z\R_DATA_TEMPR7[17] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0_DB_DETECT, 
        \Z\ACCESS_BUSY[7][0] , \Z\R_DATA_TEMPR25[44] , OR4_320_Y, 
        \Z\R_DATA_TEMPR30[15] , \Z\R_DATA_TEMPR31[15] , 
        \Z\R_DATA_TEMPR13[17] , \Z\R_DATA_TEMPR15[17] , OR4_331_Y, 
        \Z\R_DATA_TEMPR16[27] , \Z\R_DATA_TEMPR17[27] , OR4_4_Y, 
        \Z\R_DATA_TEMPR24[24] , \Z\R_DATA_TEMPR25[24] , 
        \Z\R_DATA_TEMPR26[24] , \Z\R_DATA_TEMPR27[24] , 
        \Z\R_DATA_TEMPR8[34] , \Z\R_DATA_TEMPR29[71] , 
        \Z\R_DATA_TEMPR30[71] , \Z\R_DATA_TEMPR31[71] , OR4_386_Y, 
        \Z\R_DATA_TEMPR16[19] , \Z\R_DATA_TEMPR17[19] , OR4_16_Y, 
        \Z\R_DATA_TEMPR13[1] , \Z\R_DATA_TEMPR15[1] , 
        \Z\R_DATA_TEMPR16[18] , \Z\R_DATA_TEMPR17[18] , OR4_100_Y, 
        OR4_149_Y, OR4_387_Y, OR4_145_Y, \Z\R_DATA_TEMPR13[10] , 
        \Z\R_DATA_TEMPR15[10] , \Z\R_DATA_TEMPR5[62] , 
        \Z\R_DATA_TEMPR7[62] , OR2_9_Y, OR4_484_Y, 
        \Z\R_DATA_TEMPR0[57] , \Z\R_DATA_TEMPR1[57] , 
        \Z\R_DATA_TEMPR2[57] , \Z\R_DATA_TEMPR3[57] , OR4_211_Y, 
        \Z\R_DATA_TEMPR16[7] , \Z\R_DATA_TEMPR17[7] , 
        \Z\R_DATA_TEMPR0[70] , \Z\R_DATA_TEMPR1[70] , 
        \Z\R_DATA_TEMPR2[70] , \Z\R_DATA_TEMPR3[70] , OR4_534_Y, 
        OR4_475_Y, OR4_317_Y, OR4_485_Y, OR4_82_Y, 
        \Z\R_DATA_TEMPR25[74] , OR4_466_Y, \Z\R_DATA_TEMPR8[23] , 
        OR4_152_Y, \Z\R_DATA_TEMPR12[54] , \Z\R_DATA_TEMPR15[54] , 
        OR4_521_Y, OR2_75_Y, \Z\R_DATA_TEMPR22[53] , 
        \Z\R_DATA_TEMPR23[53] , OR4_358_Y, OR4_499_Y, OR4_551_Y, 
        \Z\R_DATA_TEMPR24[35] , \Z\R_DATA_TEMPR25[35] , 
        \Z\R_DATA_TEMPR26[35] , \Z\R_DATA_TEMPR27[35] , OR2_55_Y, 
        \Z\R_DATA_TEMPR19[66] , \Z\R_DATA_TEMPR16[4] , 
        \Z\R_DATA_TEMPR17[4] , \Z\R_DATA_TEMPR25[58] , OR4_568_Y, 
        \Z\R_DATA_TEMPR4[0] , \Z\R_DATA_TEMPR6[0] , 
        \Z\R_DATA_TEMPR8[20] , \Z\R_DATA_TEMPR21[63] , OR4_174_Y, 
        \Z\R_DATA_TEMPR13[6] , \Z\R_DATA_TEMPR15[6] , OR4_292_Y, 
        \Z\R_DATA_TEMPR29[62] , \Z\R_DATA_TEMPR30[62] , 
        \Z\R_DATA_TEMPR31[62] , \Z\R_DATA_TEMPR21[72] , OR4_104_Y, 
        \Z\R_DATA_TEMPR16[26] , \Z\R_DATA_TEMPR17[26] , 
        \Z\R_DATA_TEMPR4[20] , \Z\R_DATA_TEMPR4[21] , 
        \Z\R_DATA_TEMPR4[22] , \Z\R_DATA_TEMPR4[23] , 
        \Z\R_DATA_TEMPR4[26] , \Z\R_DATA_TEMPR4[28] , 
        \Z\R_DATA_TEMPR4[29] , \Z\R_DATA_TEMPR4[30] , 
        \Z\R_DATA_TEMPR4[31] , \Z\R_DATA_TEMPR4[37] , 
        \Z\R_DATA_TEMPR4[38] , \Z\R_DATA_TEMPR4[1] , 
        \Z\R_DATA_TEMPR4[2] , \Z\R_DATA_TEMPR4[3] , 
        \Z\R_DATA_TEMPR4[4] , \Z\R_DATA_TEMPR4[5] , 
        \Z\R_DATA_TEMPR4[6] , \Z\R_DATA_TEMPR4[8] , 
        \Z\R_DATA_TEMPR4[9] , \Z\R_DATA_TEMPR4[14] , 
        \Z\R_DATA_TEMPR4[17] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0_DB_DETECT, 
        \Z\ACCESS_BUSY[4][0] , \Z\R_DATA_TEMPR6[2] , OR4_9_Y, OR2_79_Y, 
        \Z\R_DATA_TEMPR22[29] , OR2_38_Y, \Z\R_DATA_TEMPR22[47] , 
        \Z\R_DATA_TEMPR23[47] , \Z\R_DATA_TEMPR22[20] , 
        \Z\R_DATA_TEMPR22[22] , \Z\R_DATA_TEMPR22[25] , 
        \Z\R_DATA_TEMPR22[26] , \Z\R_DATA_TEMPR22[27] , 
        \Z\R_DATA_TEMPR22[28] , \Z\R_DATA_TEMPR22[31] , 
        \Z\R_DATA_TEMPR22[36] , \Z\R_DATA_TEMPR22[37] , 
        \Z\R_DATA_TEMPR22[38] , \Z\R_DATA_TEMPR22[39] , 
        \Z\R_DATA_TEMPR22[0] , \Z\R_DATA_TEMPR22[1] , 
        \Z\R_DATA_TEMPR22[2] , \Z\R_DATA_TEMPR22[3] , 
        \Z\R_DATA_TEMPR22[6] , \Z\R_DATA_TEMPR22[7] , 
        \Z\R_DATA_TEMPR22[8] , \Z\R_DATA_TEMPR22[11] , 
        \Z\R_DATA_TEMPR22[14] , \Z\R_DATA_TEMPR22[15] , 
        \Z\R_DATA_TEMPR22[17] , \Z\R_DATA_TEMPR22[19] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0_DB_DETECT, 
        \Z\ACCESS_BUSY[22][0] , \Z\R_DATA_TEMPR0[47] , 
        \Z\R_DATA_TEMPR1[47] , \Z\R_DATA_TEMPR2[47] , 
        \Z\R_DATA_TEMPR3[47] , \Z\R_DATA_TEMPR9[69] , 
        \Z\R_DATA_TEMPR10[69] , \Z\R_DATA_TEMPR11[69] , OR2_44_Y, 
        OR4_228_Y, \Z\R_DATA_TEMPR13[5] , \Z\R_DATA_TEMPR15[5] , 
        OR4_148_Y, \Z\R_DATA_TEMPR16[28] , \Z\R_DATA_TEMPR17[28] , 
        OR2_15_Y, \Z\R_DATA_TEMPR22[44] , \Z\R_DATA_TEMPR23[44] , 
        OR4_621_Y, \Z\R_DATA_TEMPR30[19] , \Z\R_DATA_TEMPR31[19] , 
        \Z\R_DATA_TEMPR13[21] , \Z\R_DATA_TEMPR15[21] , 
        \Z\R_DATA_TEMPR5[44] , \Z\R_DATA_TEMPR7[44] , OR4_653_Y, 
        \Z\R_DATA_TEMPR13[31] , \Z\R_DATA_TEMPR15[31] , 
        \Z\R_DATA_TEMPR16[30] , \Z\R_DATA_TEMPR17[30] , 
        \Z\R_DATA_TEMPR2[2] , OR4_140_Y, \Z\R_DATA_TEMPR16[6] , 
        \Z\R_DATA_TEMPR17[6] , \Z\R_DATA_TEMPR8[19] , OR4_555_Y, 
        \Z\R_DATA_TEMPR16[39] , \Z\R_DATA_TEMPR17[39] , 
        \Z\R_DATA_TEMPR6[4] , OR4_404_Y, \Z\R_DATA_TEMPR0[65] , 
        \Z\R_DATA_TEMPR1[65] , \Z\R_DATA_TEMPR2[65] , 
        \Z\R_DATA_TEMPR3[65] , OR4_164_Y, \Z\R_DATA_TEMPR24[23] , 
        \Z\R_DATA_TEMPR25[23] , \Z\R_DATA_TEMPR26[23] , 
        \Z\R_DATA_TEMPR27[23] , OR4_235_Y, OR4_180_Y, 
        \Z\R_DATA_TEMPR8[21] , \Z\R_DATA_TEMPR8[24] , 
        \Z\R_DATA_TEMPR8[28] , \Z\R_DATA_TEMPR8[29] , 
        \Z\R_DATA_TEMPR8[30] , \Z\R_DATA_TEMPR8[31] , 
        \Z\R_DATA_TEMPR8[32] , \Z\R_DATA_TEMPR8[37] , 
        \Z\R_DATA_TEMPR8[38] , \Z\R_DATA_TEMPR8[3] , 
        \Z\R_DATA_TEMPR8[4] , \Z\R_DATA_TEMPR8[5] , 
        \Z\R_DATA_TEMPR8[6] , \Z\R_DATA_TEMPR8[8] , 
        \Z\R_DATA_TEMPR8[9] , \Z\R_DATA_TEMPR8[10] , 
        \Z\R_DATA_TEMPR8[11] , \Z\R_DATA_TEMPR8[14] , 
        \Z\R_DATA_TEMPR8[15] , \Z\R_DATA_TEMPR8[17] , 
        \Z\R_DATA_TEMPR8[18] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0_DB_DETECT, 
        \Z\ACCESS_BUSY[8][0] , OR4_640_Y, \Z\R_DATA_TEMPR9[51] , 
        \Z\R_DATA_TEMPR10[51] , \Z\R_DATA_TEMPR11[51] , OR4_28_Y, 
        \Z\R_DATA_TEMPR25[65] , OR4_87_Y, OR4_433_Y, OR4_692_Y, 
        OR4_298_Y, \Z\R_DATA_TEMPR29[75] , \Z\R_DATA_TEMPR30[75] , 
        \Z\R_DATA_TEMPR31[75] , OR4_427_Y, \Z\R_DATA_TEMPR16[1] , 
        \Z\R_DATA_TEMPR17[1] , \Z\R_DATA_TEMPR6[17] , OR4_187_Y, 
        OR2_32_Y, OR4_493_Y, \Z\R_DATA_TEMPR25[53] , OR4_488_Y, 
        OR4_365_Y, \Z\R_DATA_TEMPR2[20] , OR4_216_Y, 
        \Z\R_DATA_TEMPR0[52] , \Z\R_DATA_TEMPR1[52] , 
        \Z\R_DATA_TEMPR2[52] , \Z\R_DATA_TEMPR3[52] , OR4_405_Y, 
        \Z\R_DATA_TEMPR2[28] , \Z\R_DATA_TEMPR5[40] , 
        \Z\R_DATA_TEMPR7[40] , OR4_619_Y, \Z\R_DATA_TEMPR9[59] , 
        \Z\R_DATA_TEMPR10[59] , \Z\R_DATA_TEMPR11[59] , OR4_645_Y, 
        \Z\R_DATA_TEMPR13[16] , \Z\R_DATA_TEMPR15[16] , 
        \Z\R_DATA_TEMPR19[60] , \Z\R_DATA_TEMPR19[61] , 
        \Z\R_DATA_TEMPR19[64] , \Z\R_DATA_TEMPR19[65] , 
        \Z\R_DATA_TEMPR19[70] , \Z\R_DATA_TEMPR19[71] , 
        \Z\R_DATA_TEMPR19[72] , \Z\R_DATA_TEMPR19[73] , 
        \Z\R_DATA_TEMPR19[75] , \Z\R_DATA_TEMPR19[76] , 
        \Z\R_DATA_TEMPR19[77] , \Z\R_DATA_TEMPR19[78] , 
        \Z\R_DATA_TEMPR19[79] , \Z\R_DATA_TEMPR19[40] , 
        \Z\R_DATA_TEMPR19[41] , \Z\R_DATA_TEMPR19[45] , 
        \Z\R_DATA_TEMPR19[51] , \Z\R_DATA_TEMPR19[54] , 
        \Z\R_DATA_TEMPR19[56] , \Z\R_DATA_TEMPR19[58] , 
        \Z\R_DATA_TEMPR19[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C1_DB_DETECT, 
        \Z\ACCESS_BUSY[19][1] , OR4_45_Y, OR4_295_Y, 
        \Z\R_DATA_TEMPR9[64] , \Z\R_DATA_TEMPR10[64] , 
        \Z\R_DATA_TEMPR11[64] , \Z\R_DATA_TEMPR30[33] , 
        \Z\R_DATA_TEMPR31[33] , \Z\R_DATA_TEMPR31[61] , 
        \Z\R_DATA_TEMPR31[63] , \Z\R_DATA_TEMPR31[66] , 
        \Z\R_DATA_TEMPR31[67] , \Z\R_DATA_TEMPR31[68] , 
        \Z\R_DATA_TEMPR31[69] , \Z\R_DATA_TEMPR31[72] , 
        \Z\R_DATA_TEMPR31[73] , \Z\R_DATA_TEMPR31[74] , 
        \Z\R_DATA_TEMPR31[76] , \Z\R_DATA_TEMPR31[77] , 
        \Z\R_DATA_TEMPR31[41] , \Z\R_DATA_TEMPR31[42] , 
        \Z\R_DATA_TEMPR31[45] , \Z\R_DATA_TEMPR31[48] , 
        \Z\R_DATA_TEMPR31[49] , \Z\R_DATA_TEMPR31[50] , 
        \Z\R_DATA_TEMPR31[52] , \Z\R_DATA_TEMPR31[54] , 
        \Z\R_DATA_TEMPR31[57] , \Z\R_DATA_TEMPR31[58] , 
        \Z\R_DATA_TEMPR31[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C1_DB_DETECT, 
        \Z\ACCESS_BUSY[31][1] , \Z\R_DATA_TEMPR24[21] , 
        \Z\R_DATA_TEMPR24[25] , \Z\R_DATA_TEMPR24[26] , 
        \Z\R_DATA_TEMPR24[29] , \Z\R_DATA_TEMPR24[30] , 
        \Z\R_DATA_TEMPR24[34] , \Z\R_DATA_TEMPR24[39] , 
        \Z\R_DATA_TEMPR24[0] , \Z\R_DATA_TEMPR24[2] , 
        \Z\R_DATA_TEMPR24[5] , \Z\R_DATA_TEMPR24[6] , 
        \Z\R_DATA_TEMPR24[7] , \Z\R_DATA_TEMPR24[8] , 
        \Z\R_DATA_TEMPR24[9] , \Z\R_DATA_TEMPR24[11] , 
        \Z\R_DATA_TEMPR24[12] , \Z\R_DATA_TEMPR24[13] , 
        \Z\R_DATA_TEMPR24[14] , \Z\R_DATA_TEMPR24[15] , 
        \Z\R_DATA_TEMPR24[16] , \Z\R_DATA_TEMPR24[18] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0_DB_DETECT, 
        \Z\ACCESS_BUSY[24][0] , \Z\R_DATA_TEMPR25[66] , OR4_517_Y, 
        \Z\R_DATA_TEMPR0[51] , \Z\R_DATA_TEMPR1[51] , 
        \Z\R_DATA_TEMPR2[51] , \Z\R_DATA_TEMPR3[51] , 
        \Z\R_DATA_TEMPR25[61] , OR4_421_Y, OR4_241_Y, OR4_294_Y, 
        OR4_464_Y, \Z\R_DATA_TEMPR0[61] , \Z\R_DATA_TEMPR1[61] , 
        \Z\R_DATA_TEMPR2[61] , \Z\R_DATA_TEMPR3[61] , 
        \Z\R_DATA_TEMPR21[78] , \Z\R_DATA_TEMPR29[58] , 
        \Z\R_DATA_TEMPR30[58] , OR4_497_Y, \Z\R_DATA_TEMPR5[78] , 
        \Z\R_DATA_TEMPR7[78] , OR2_65_Y, \Z\R_DATA_TEMPR0[77] , 
        \Z\R_DATA_TEMPR1[77] , \Z\R_DATA_TEMPR2[77] , 
        \Z\R_DATA_TEMPR3[77] , \Z\R_DATA_TEMPR13[36] , 
        \Z\R_DATA_TEMPR15[36] , \Z\R_DATA_TEMPR21[69] , OR4_236_Y, 
        \Z\R_DATA_TEMPR25[13] , \Z\R_DATA_TEMPR26[13] , 
        \Z\R_DATA_TEMPR27[13] , OR4_345_Y, \Z\R_DATA_TEMPR16[31] , 
        \Z\R_DATA_TEMPR17[31] , \Z\R_DATA_TEMPR6[9] , OR4_11_Y, 
        \Z\R_DATA_TEMPR6[1] , \Z\R_DATA_TEMPR23[64] , 
        \Z\R_DATA_TEMPR23[68] , \Z\R_DATA_TEMPR23[73] , 
        \Z\R_DATA_TEMPR23[74] , \Z\R_DATA_TEMPR23[76] , 
        \Z\R_DATA_TEMPR23[77] , \Z\R_DATA_TEMPR23[79] , 
        \Z\R_DATA_TEMPR23[40] , \Z\R_DATA_TEMPR23[41] , 
        \Z\R_DATA_TEMPR23[42] , \Z\R_DATA_TEMPR23[43] , 
        \Z\R_DATA_TEMPR23[45] , \Z\R_DATA_TEMPR23[48] , 
        \Z\R_DATA_TEMPR23[49] , \Z\R_DATA_TEMPR23[50] , 
        \Z\R_DATA_TEMPR23[52] , \Z\R_DATA_TEMPR23[54] , 
        \Z\R_DATA_TEMPR23[55] , \Z\R_DATA_TEMPR23[56] , 
        \Z\R_DATA_TEMPR23[58] , \Z\R_DATA_TEMPR23[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C1_DB_DETECT, 
        \Z\ACCESS_BUSY[23][1] , \Z\R_DATA_TEMPR9[53] , 
        \Z\R_DATA_TEMPR10[53] , \Z\R_DATA_TEMPR11[53] , 
        \Z\R_DATA_TEMPR30[2] , \Z\R_DATA_TEMPR31[2] , OR4_312_Y, 
        \Z\R_DATA_TEMPR30[4] , \Z\R_DATA_TEMPR31[4] , 
        \Z\R_DATA_TEMPR9[58] , \Z\R_DATA_TEMPR10[58] , 
        \Z\R_DATA_TEMPR11[58] , \Z\R_DATA_TEMPR16[16] , 
        \Z\R_DATA_TEMPR17[16] , \Z\R_DATA_TEMPR17[21] , 
        \Z\R_DATA_TEMPR17[22] , \Z\R_DATA_TEMPR17[32] , 
        \Z\R_DATA_TEMPR17[33] , \Z\R_DATA_TEMPR17[34] , 
        \Z\R_DATA_TEMPR17[38] , \Z\R_DATA_TEMPR17[0] , 
        \Z\R_DATA_TEMPR17[3] , \Z\R_DATA_TEMPR17[5] , 
        \Z\R_DATA_TEMPR17[8] , \Z\R_DATA_TEMPR17[9] , 
        \Z\R_DATA_TEMPR17[10] , \Z\R_DATA_TEMPR17[11] , 
        \Z\R_DATA_TEMPR17[12] , \Z\R_DATA_TEMPR17[13] , 
        \Z\R_DATA_TEMPR17[14] , \Z\R_DATA_TEMPR17[15] , 
        \Z\R_DATA_TEMPR17[17] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0_DB_DETECT, 
        \Z\ACCESS_BUSY[17][0] , OR2_42_Y, OR4_537_Y, 
        \Z\R_DATA_TEMPR5[68] , \Z\R_DATA_TEMPR7[68] , OR4_590_Y, 
        OR4_128_Y, \Z\R_DATA_TEMPR16[22] , \Z\R_DATA_TEMPR15[20] , 
        \Z\R_DATA_TEMPR15[22] , \Z\R_DATA_TEMPR15[23] , 
        \Z\R_DATA_TEMPR15[24] , \Z\R_DATA_TEMPR15[28] , 
        \Z\R_DATA_TEMPR15[29] , \Z\R_DATA_TEMPR15[32] , 
        \Z\R_DATA_TEMPR15[33] , \Z\R_DATA_TEMPR15[35] , 
        \Z\R_DATA_TEMPR15[39] , \Z\R_DATA_TEMPR15[0] , 
        \Z\R_DATA_TEMPR15[2] , \Z\R_DATA_TEMPR15[3] , 
        \Z\R_DATA_TEMPR15[4] , \Z\R_DATA_TEMPR15[9] , 
        \Z\R_DATA_TEMPR15[11] , \Z\R_DATA_TEMPR15[14] , 
        \Z\R_DATA_TEMPR15[15] , \Z\R_DATA_TEMPR15[18] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0_DB_DETECT, 
        \Z\ACCESS_BUSY[15][0] , \Z\R_DATA_TEMPR13[20] , 
        \Z\R_DATA_TEMPR25[6] , \Z\R_DATA_TEMPR26[6] , 
        \Z\R_DATA_TEMPR27[6] , OR2_58_Y, \Z\R_DATA_TEMPR13[18] , 
        OR4_673_Y, OR4_68_Y, OR4_416_Y, \Z\R_DATA_TEMPR30[21] , 
        \Z\R_DATA_TEMPR31[21] , OR2_39_Y, \Z\R_DATA_TEMPR6[29] , 
        OR4_707_Y, \Z\R_DATA_TEMPR29[45] , \Z\R_DATA_TEMPR30[45] , 
        OR2_69_Y, OR4_698_Y, OR4_26_Y, OR2_2_Y, \Z\R_DATA_TEMPR21[52] , 
        OR4_51_Y, \Z\R_DATA_TEMPR9[52] , \Z\R_DATA_TEMPR10[52] , 
        \Z\R_DATA_TEMPR11[52] , \Z\R_DATA_TEMPR29[41] , 
        \Z\R_DATA_TEMPR30[41] , OR4_327_Y, \Z\R_DATA_TEMPR6[6] , 
        \Z\R_DATA_TEMPR0[62] , \Z\R_DATA_TEMPR1[62] , 
        \Z\R_DATA_TEMPR2[62] , \Z\R_DATA_TEMPR3[62] , OR4_518_Y, 
        OR4_247_Y, OR4_106_Y, OR4_13_Y, \Z\R_DATA_TEMPR29[48] , 
        \Z\R_DATA_TEMPR30[48] , OR4_332_Y, \Z\R_DATA_TEMPR30[36] , 
        \Z\R_DATA_TEMPR31[36] , OR4_183_Y, OR4_305_Y, OR4_159_Y, 
        OR4_620_Y, \Z\R_DATA_TEMPR12[43] , \Z\R_DATA_TEMPR15[43] , 
        OR4_647_Y, OR2_49_Y, OR4_258_Y, \Z\R_DATA_TEMPR22[48] , 
        \Z\R_DATA_TEMPR5[50] , \Z\R_DATA_TEMPR7[50] , OR4_279_Y, 
        OR4_89_Y, OR4_453_Y, \Z\R_DATA_TEMPR6[3] , OR4_436_Y, 
        OR4_658_Y, OR4_435_Y, OR4_420_Y, OR2_66_Y, 
        \Z\R_DATA_TEMPR22[56] , \Z\R_DATA_TEMPR2[23] , 
        \Z\R_DATA_TEMPR2[24] , \Z\R_DATA_TEMPR2[27] , 
        \Z\R_DATA_TEMPR2[29] , \Z\R_DATA_TEMPR2[30] , 
        \Z\R_DATA_TEMPR2[31] , \Z\R_DATA_TEMPR2[35] , 
        \Z\R_DATA_TEMPR2[36] , \Z\R_DATA_TEMPR2[39] , 
        \Z\R_DATA_TEMPR2[1] , \Z\R_DATA_TEMPR2[3] , 
        \Z\R_DATA_TEMPR2[6] , \Z\R_DATA_TEMPR2[7] , 
        \Z\R_DATA_TEMPR2[8] , \Z\R_DATA_TEMPR2[9] , 
        \Z\R_DATA_TEMPR2[11] , \Z\R_DATA_TEMPR2[12] , 
        \Z\R_DATA_TEMPR2[15] , \Z\R_DATA_TEMPR2[17] , 
        \Z\R_DATA_TEMPR2[18] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0_DB_DETECT, 
        \Z\ACCESS_BUSY[2][0] , \Z\R_DATA_TEMPR15[67] , 
        \Z\R_DATA_TEMPR15[69] , \Z\R_DATA_TEMPR15[70] , 
        \Z\R_DATA_TEMPR15[72] , \Z\R_DATA_TEMPR15[73] , 
        \Z\R_DATA_TEMPR15[74] , \Z\R_DATA_TEMPR15[75] , 
        \Z\R_DATA_TEMPR15[76] , \Z\R_DATA_TEMPR15[77] , 
        \Z\R_DATA_TEMPR15[40] , \Z\R_DATA_TEMPR15[41] , 
        \Z\R_DATA_TEMPR15[45] , \Z\R_DATA_TEMPR15[46] , 
        \Z\R_DATA_TEMPR15[47] , \Z\R_DATA_TEMPR15[50] , 
        \Z\R_DATA_TEMPR15[51] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C1_DB_DETECT, 
        \Z\ACCESS_BUSY[15][1] , OR4_516_Y, OR4_300_Y, OR4_349_Y, 
        \Z\R_DATA_TEMPR16[12] , \Z\R_DATA_TEMPR0[60] , 
        \Z\R_DATA_TEMPR0[66] , \Z\R_DATA_TEMPR0[68] , 
        \Z\R_DATA_TEMPR0[72] , \Z\R_DATA_TEMPR0[74] , 
        \Z\R_DATA_TEMPR0[79] , \Z\R_DATA_TEMPR0[40] , 
        \Z\R_DATA_TEMPR0[42] , \Z\R_DATA_TEMPR0[43] , 
        \Z\R_DATA_TEMPR0[44] , \Z\R_DATA_TEMPR0[45] , 
        \Z\R_DATA_TEMPR0[49] , \Z\R_DATA_TEMPR0[53] , 
        \Z\R_DATA_TEMPR0[54] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C1_DB_DETECT, 
        \Z\ACCESS_BUSY[0][1] , OR4_683_Y, \Z\R_DATA_TEMPR1[68] , 
        \Z\R_DATA_TEMPR2[68] , \Z\R_DATA_TEMPR3[68] , OR4_53_Y, 
        \Z\R_DATA_TEMPR6[37] , \Z\R_DATA_TEMPR30[20] , 
        \Z\R_DATA_TEMPR31[20] , OR4_538_Y, OR4_625_Y, 
        \Z\R_DATA_TEMPR5[52] , \Z\R_DATA_TEMPR7[52] , OR4_397_Y, 
        \Z\R_DATA_TEMPR16[17] , \Z\R_DATA_TEMPR30[32] , 
        \Z\R_DATA_TEMPR31[32] , \Z\R_DATA_TEMPR13[29] , OR4_711_Y, 
        OR4_88_Y, OR4_628_Y, OR4_603_Y, \Z\R_DATA_TEMPR25[21] , 
        \Z\R_DATA_TEMPR26[21] , \Z\R_DATA_TEMPR27[21] , OR4_277_Y, 
        OR4_172_Y, \Z\R_DATA_TEMPR13[28] , OR4_675_Y, OR4_310_Y, 
        \Z\R_DATA_TEMPR25[5] , \Z\R_DATA_TEMPR26[5] , 
        \Z\R_DATA_TEMPR27[5] , OR4_218_Y, OR4_42_Y, OR4_714_Y, 
        OR2_57_Y, \Z\R_DATA_TEMPR21[73] , OR4_155_Y, 
        \Z\R_DATA_TEMPR5[55] , \Z\R_DATA_TEMPR7[55] , 
        \Z\R_DATA_TEMPR5[46] , \Z\R_DATA_TEMPR7[46] , 
        \Z\R_DATA_TEMPR21[60] , OR4_325_Y, \Z\R_DATA_TEMPR1[43] , 
        \Z\R_DATA_TEMPR2[43] , \Z\R_DATA_TEMPR3[43] , OR4_377_Y, 
        OR2_37_Y, OR4_62_Y, OR4_695_Y, \Z\R_DATA_TEMPR16[15] , 
        OR4_269_Y, \Z\R_DATA_TEMPR12[75] , OR4_156_Y, OR4_49_Y, 
        OR4_448_Y, \Z\R_DATA_TEMPR30[16] , \Z\R_DATA_TEMPR31[16] , 
        OR4_434_Y, OR4_219_Y, \Z\R_DATA_TEMPR30[14] , 
        \Z\R_DATA_TEMPR31[14] , \Z\R_DATA_TEMPR6[8] , OR4_224_Y, 
        OR4_103_Y, \Z\R_DATA_TEMPR29[69] , \Z\R_DATA_TEMPR30[69] , 
        OR2_35_Y, \Z\R_DATA_TEMPR12[69] , OR4_316_Y, OR4_328_Y, 
        \Z\R_DATA_TEMPR16[21] , \Z\R_DATA_TEMPR16[32] , 
        \Z\R_DATA_TEMPR16[33] , \Z\R_DATA_TEMPR16[34] , 
        \Z\R_DATA_TEMPR16[38] , \Z\R_DATA_TEMPR16[0] , 
        \Z\R_DATA_TEMPR16[3] , \Z\R_DATA_TEMPR16[5] , 
        \Z\R_DATA_TEMPR16[8] , \Z\R_DATA_TEMPR16[9] , 
        \Z\R_DATA_TEMPR16[10] , \Z\R_DATA_TEMPR16[11] , 
        \Z\R_DATA_TEMPR16[13] , \Z\R_DATA_TEMPR16[14] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0_DB_DETECT, 
        \Z\ACCESS_BUSY[16][0] , OR4_282_Y, OR4_565_Y, OR4_663_Y, 
        \Z\R_DATA_TEMPR12[47] , \Z\R_DATA_TEMPR30[61] , 
        \Z\R_DATA_TEMPR30[63] , \Z\R_DATA_TEMPR30[66] , 
        \Z\R_DATA_TEMPR30[67] , \Z\R_DATA_TEMPR30[68] , 
        \Z\R_DATA_TEMPR30[72] , \Z\R_DATA_TEMPR30[73] , 
        \Z\R_DATA_TEMPR30[74] , \Z\R_DATA_TEMPR30[76] , 
        \Z\R_DATA_TEMPR30[77] , \Z\R_DATA_TEMPR30[42] , 
        \Z\R_DATA_TEMPR30[49] , \Z\R_DATA_TEMPR30[50] , 
        \Z\R_DATA_TEMPR30[52] , \Z\R_DATA_TEMPR30[54] , 
        \Z\R_DATA_TEMPR30[57] , \Z\R_DATA_TEMPR30[59] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C1_DB_DETECT, 
        \Z\ACCESS_BUSY[30][1] , \Z\R_DATA_TEMPR29[74] , OR4_127_Y, 
        \Z\R_DATA_TEMPR9[65] , \Z\R_DATA_TEMPR10[65] , 
        \Z\R_DATA_TEMPR11[65] , \Z\R_DATA_TEMPR12[50] , OR4_395_Y, 
        \Z\R_DATA_TEMPR25[49] , \Z\R_DATA_TEMPR12[73] , OR4_69_Y, 
        \Z\R_DATA_TEMPR30[12] , \Z\R_DATA_TEMPR31[12] , 
        \Z\R_DATA_TEMPR25[43] , \Z\R_DATA_TEMPR21[57] , OR4_575_Y, 
        \Z\R_DATA_TEMPR6[5] , OR4_581_Y, \Z\R_DATA_TEMPR12[74] , 
        OR4_398_Y, OR4_158_Y, \Z\R_DATA_TEMPR5[57] , 
        \Z\R_DATA_TEMPR7[57] , OR4_146_Y, OR4_85_Y, 
        \Z\R_DATA_TEMPR13[39] , OR4_505_Y, \Z\R_DATA_TEMPR25[75] , 
        OR4_449_Y, \Z\R_DATA_TEMPR13[35] , \Z\R_DATA_TEMPR29[57] , 
        OR4_415_Y, OR4_336_Y, OR4_655_Y, \Z\R_DATA_TEMPR22[59] , 
        OR4_343_Y, OR4_163_Y, \Z\R_DATA_TEMPR29[59] , OR4_357_Y, 
        OR4_197_Y, \Z\R_DATA_TEMPR13[23] , OR4_37_Y, OR4_703_Y, 
        OR4_549_Y, \Z\R_DATA_TEMPR6[22] , \Z\R_DATA_TEMPR9[60] , 
        \Z\R_DATA_TEMPR9[62] , \Z\R_DATA_TEMPR9[63] , 
        \Z\R_DATA_TEMPR9[66] , \Z\R_DATA_TEMPR9[67] , 
        \Z\R_DATA_TEMPR9[68] , \Z\R_DATA_TEMPR9[73] , 
        \Z\R_DATA_TEMPR9[74] , \Z\R_DATA_TEMPR9[76] , 
        \Z\R_DATA_TEMPR9[40] , \Z\R_DATA_TEMPR9[42] , 
        \Z\R_DATA_TEMPR9[43] , \Z\R_DATA_TEMPR9[44] , 
        \Z\R_DATA_TEMPR9[46] , \Z\R_DATA_TEMPR9[55] , 
        \Z\R_DATA_TEMPR9[57] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C1_DB_DETECT, 
        \Z\ACCESS_BUSY[9][1] , OR4_627_Y, OR2_8_Y, 
        \Z\R_DATA_TEMPR22[45] , OR4_650_Y, \Z\R_DATA_TEMPR29[54] , 
        OR4_30_Y, \Z\R_DATA_TEMPR1[60] , \Z\R_DATA_TEMPR2[60] , 
        \Z\R_DATA_TEMPR3[60] , OR4_708_Y, OR4_324_Y, 
        \Z\R_DATA_TEMPR29[61] , \Z\R_DATA_TEMPR29[63] , 
        \Z\R_DATA_TEMPR29[66] , \Z\R_DATA_TEMPR29[67] , 
        \Z\R_DATA_TEMPR29[68] , \Z\R_DATA_TEMPR29[72] , 
        \Z\R_DATA_TEMPR29[73] , \Z\R_DATA_TEMPR29[76] , 
        \Z\R_DATA_TEMPR29[77] , \Z\R_DATA_TEMPR29[42] , 
        \Z\R_DATA_TEMPR29[49] , \Z\R_DATA_TEMPR29[50] , 
        \Z\R_DATA_TEMPR29[52] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C1_DB_DETECT, 
        \Z\ACCESS_BUSY[29][1] , OR4_370_Y, \Z\R_DATA_TEMPR12[45] , 
        OR4_681_Y, \Z\R_DATA_TEMPR25[29] , \Z\R_DATA_TEMPR26[29] , 
        \Z\R_DATA_TEMPR27[29] , OR4_483_Y, OR4_540_Y, 
        \Z\R_DATA_TEMPR6[31] , \Z\R_DATA_TEMPR22[50] , 
        \Z\R_DATA_TEMPR25[63] , \Z\R_DATA_TEMPR6[30] , OR4_44_Y, 
        \Z\R_DATA_TEMPR22[52] , \Z\R_DATA_TEMPR1[45] , 
        \Z\R_DATA_TEMPR2[45] , \Z\R_DATA_TEMPR3[45] , OR4_272_Y, 
        \Z\R_DATA_TEMPR25[18] , \Z\R_DATA_TEMPR26[18] , 
        \Z\R_DATA_TEMPR27[18] , OR4_253_Y, \Z\R_DATA_TEMPR25[39] , 
        \Z\R_DATA_TEMPR26[39] , \Z\R_DATA_TEMPR27[39] , OR4_479_Y, 
        \Z\R_DATA_TEMPR25[16] , \Z\R_DATA_TEMPR26[16] , 
        \Z\R_DATA_TEMPR27[16] , OR4_21_Y, \Z\R_DATA_TEMPR10[63] , 
        \Z\R_DATA_TEMPR11[63] , \Z\R_DATA_TEMPR27[25] , 
        \Z\R_DATA_TEMPR27[26] , \Z\R_DATA_TEMPR27[30] , 
        \Z\R_DATA_TEMPR27[34] , \Z\R_DATA_TEMPR27[0] , 
        \Z\R_DATA_TEMPR27[2] , \Z\R_DATA_TEMPR27[7] , 
        \Z\R_DATA_TEMPR27[8] , \Z\R_DATA_TEMPR27[9] , 
        \Z\R_DATA_TEMPR27[11] , \Z\R_DATA_TEMPR27[12] , 
        \Z\R_DATA_TEMPR27[14] , \Z\R_DATA_TEMPR27[15] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0_DB_DETECT, 
        \Z\ACCESS_BUSY[27][0] , OR2_47_Y, \Z\R_DATA_TEMPR25[79] , 
        \Z\R_DATA_TEMPR10[76] , \Z\R_DATA_TEMPR11[76] , OR4_36_Y, 
        \Z\R_DATA_TEMPR10[60] , \Z\R_DATA_TEMPR11[60] , OR4_607_Y, 
        OR4_440_Y, OR4_278_Y, \Z\R_DATA_TEMPR25[25] , 
        \Z\R_DATA_TEMPR25[26] , \Z\R_DATA_TEMPR25[30] , 
        \Z\R_DATA_TEMPR25[34] , \Z\R_DATA_TEMPR25[0] , 
        \Z\R_DATA_TEMPR25[2] , \Z\R_DATA_TEMPR25[7] , 
        \Z\R_DATA_TEMPR25[8] , \Z\R_DATA_TEMPR25[9] , 
        \Z\R_DATA_TEMPR25[11] , \Z\R_DATA_TEMPR25[12] , 
        \Z\R_DATA_TEMPR25[14] , \Z\R_DATA_TEMPR25[15] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0_DB_DETECT, 
        \Z\ACCESS_BUSY[25][0] , OR4_185_Y, \Z\R_DATA_TEMPR10[43] , 
        \Z\R_DATA_TEMPR11[43] , OR4_344_Y, OR4_94_Y, 
        \Z\R_DATA_TEMPR5[65] , \Z\R_DATA_TEMPR7[65] , OR4_126_Y, 
        OR4_262_Y, OR4_429_Y, \Z\R_DATA_TEMPR10[57] , 
        \Z\R_DATA_TEMPR11[57] , OR4_254_Y, \Z\R_DATA_TEMPR13[3] , 
        \Z\R_DATA_TEMPR1[40] , \Z\R_DATA_TEMPR2[40] , 
        \Z\R_DATA_TEMPR3[40] , OR4_23_Y, \Z\R_DATA_TEMPR5[41] , 
        \Z\R_DATA_TEMPR7[41] , OR4_422_Y, OR4_696_Y, OR4_605_Y, 
        \Z\R_DATA_TEMPR21[47] , OR4_671_Y, \Z\R_DATA_TEMPR25[52] , 
        \Z\R_DATA_TEMPR22[77] , OR4_66_Y, OR4_191_Y, OR4_83_Y, 
        OR4_482_Y, OR4_580_Y, \Z\R_DATA_TEMPR25[70] , 
        \Z\R_DATA_TEMPR30[13] , \Z\R_DATA_TEMPR31[13] , OR4_208_Y, 
        \Z\R_DATA_TEMPR30[37] , \Z\R_DATA_TEMPR31[37] , OR2_68_Y, 
        \Z\R_DATA_TEMPR30[5] , \Z\R_DATA_TEMPR31[5] , 
        \Z\R_DATA_TEMPR22[40] , OR4_561_Y, \Z\R_DATA_TEMPR30[29] , 
        \Z\R_DATA_TEMPR31[29] , \Z\R_DATA_TEMPR5[60] , 
        \Z\R_DATA_TEMPR5[61] , \Z\R_DATA_TEMPR5[63] , 
        \Z\R_DATA_TEMPR5[66] , \Z\R_DATA_TEMPR5[67] , 
        \Z\R_DATA_TEMPR5[69] , \Z\R_DATA_TEMPR5[79] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C1_DB_DETECT, 
        \Z\ACCESS_BUSY[5][1] , \Z\R_DATA_TEMPR13[9] , 
        \Z\R_DATA_TEMPR26[12] , \Z\R_DATA_TEMPR25[67] , 
        \Z\R_DATA_TEMPR25[68] , \Z\R_DATA_TEMPR25[69] , 
        \Z\R_DATA_TEMPR25[77] , \Z\R_DATA_TEMPR25[42] , 
        \Z\R_DATA_TEMPR25[47] , \Z\R_DATA_TEMPR25[54] , 
        \Z\R_DATA_TEMPR25[57] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C1_DB_DETECT, 
        \Z\ACCESS_BUSY[25][1] , OR4_670_Y, \Z\R_DATA_TEMPR26[8] , 
        OR2_48_Y, \Z\R_DATA_TEMPR21[49] , OR4_112_Y, OR4_196_Y, 
        \Z\R_DATA_TEMPR10[55] , \Z\R_DATA_TEMPR11[55] , 
        \Z\R_DATA_TEMPR1[66] , \Z\R_DATA_TEMPR2[66] , 
        \Z\R_DATA_TEMPR3[66] , \Z\R_DATA_TEMPR26[2] , 
        \Z\R_DATA_TEMPR22[55] , OR4_492_Y, \Z\R_DATA_TEMPR1[79] , 
        \Z\R_DATA_TEMPR2[79] , \Z\R_DATA_TEMPR3[79] , OR4_477_Y, 
        \Z\R_DATA_TEMPR6[23] , OR4_529_Y, \Z\R_DATA_TEMPR26[30] , 
        OR2_33_Y, \Z\R_DATA_TEMPR22[79] , OR4_685_Y, OR4_175_Y, 
        \Z\R_DATA_TEMPR6[26] , OR4_268_Y, \Z\R_DATA_TEMPR6[28] , 
        OR4_631_Y, OR4_661_Y, \Z\R_DATA_TEMPR13[4] , 
        \Z\R_DATA_TEMPR11[62] , \Z\R_DATA_TEMPR11[66] , 
        \Z\R_DATA_TEMPR11[67] , \Z\R_DATA_TEMPR11[68] , 
        \Z\R_DATA_TEMPR11[73] , \Z\R_DATA_TEMPR11[74] , 
        \Z\R_DATA_TEMPR11[40] , \Z\R_DATA_TEMPR11[42] , 
        \Z\R_DATA_TEMPR11[44] , \Z\R_DATA_TEMPR11[46] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C1_DB_DETECT, 
        \Z\ACCESS_BUSY[11][1] , OR4_7_Y, \Z\R_DATA_TEMPR7[79] , 
        OR4_132_Y, \Z\R_DATA_TEMPR1[72] , \Z\R_DATA_TEMPR1[74] , 
        \Z\R_DATA_TEMPR1[42] , \Z\R_DATA_TEMPR1[44] , 
        \Z\R_DATA_TEMPR1[49] , \Z\R_DATA_TEMPR1[53] , 
        \Z\R_DATA_TEMPR1[54] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C1_DB_DETECT, 
        \Z\ACCESS_BUSY[1][1] , OR4_99_Y, \Z\R_DATA_TEMPR3[72] , 
        \Z\R_DATA_TEMPR3[74] , \Z\R_DATA_TEMPR3[42] , 
        \Z\R_DATA_TEMPR3[44] , \Z\R_DATA_TEMPR3[49] , 
        \Z\R_DATA_TEMPR3[53] , \Z\R_DATA_TEMPR3[54] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C1_DB_DETECT, 
        \Z\ACCESS_BUSY[3][1] , \Z\R_DATA_TEMPR21[65] , 
        \Z\R_DATA_TEMPR30[25] , \Z\R_DATA_TEMPR30[27] , 
        \Z\R_DATA_TEMPR30[30] , \Z\R_DATA_TEMPR30[31] , 
        \Z\R_DATA_TEMPR30[38] , \Z\R_DATA_TEMPR30[1] , 
        \Z\R_DATA_TEMPR30[6] , \Z\R_DATA_TEMPR30[7] , 
        \Z\R_DATA_TEMPR30[8] , \Z\R_DATA_TEMPR30[11] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0_DB_DETECT, 
        \Z\ACCESS_BUSY[30][0] , \Z\R_DATA_TEMPR7[61] , OR4_702_Y, 
        OR4_265_Y, OR4_642_Y, \Z\R_DATA_TEMPR26[25] , 
        \Z\R_DATA_TEMPR26[26] , \Z\R_DATA_TEMPR26[34] , 
        \Z\R_DATA_TEMPR26[0] , \Z\R_DATA_TEMPR26[7] , 
        \Z\R_DATA_TEMPR26[9] , \Z\R_DATA_TEMPR26[11] , 
        \Z\R_DATA_TEMPR26[14] , \Z\R_DATA_TEMPR26[15] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0_DB_DETECT, 
        \Z\ACCESS_BUSY[26][0] , \Z\R_DATA_TEMPR12[76] , OR2_74_Y, 
        OR2_60_Y, \Z\R_DATA_TEMPR21[64] , OR4_648_Y, 
        \Z\R_DATA_TEMPR31[31] , OR4_176_Y, OR4_92_Y, 
        \Z\R_DATA_TEMPR10[73] , OR2_19_Y, \Z\R_DATA_TEMPR22[58] , 
        OR4_491_Y, \Z\R_DATA_TEMPR13[11] , \Z\R_DATA_TEMPR10[42] , 
        OR4_264_Y, OR4_151_Y, OR2_40_Y, \Z\R_DATA_TEMPR10[66] , 
        \Z\R_DATA_TEMPR12[67] , \Z\R_DATA_TEMPR12[70] , 
        \Z\R_DATA_TEMPR12[72] , \Z\R_DATA_TEMPR12[77] , 
        \Z\R_DATA_TEMPR12[40] , \Z\R_DATA_TEMPR12[41] , 
        \Z\R_DATA_TEMPR12[46] , \Z\R_DATA_TEMPR12[51] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C1_DB_DETECT, 
        \Z\ACCESS_BUSY[12][1] , OR4_413_Y, \Z\R_DATA_TEMPR13[22] , 
        OR2_46_Y, OR4_243_Y, \Z\R_DATA_TEMPR10[67] , OR4_170_Y, 
        OR4_115_Y, OR4_31_Y, \Z\R_DATA_TEMPR7[63] , 
        \Z\R_DATA_TEMPR2[72] , \Z\R_DATA_TEMPR22[54] , OR4_535_Y, 
        \Z\R_DATA_TEMPR22[42] , OR4_459_Y, \Z\R_DATA_TEMPR21[56] , 
        \Z\R_DATA_TEMPR13[32] , \Z\R_DATA_TEMPR13[15] , OR4_600_Y, 
        \Z\R_DATA_TEMPR7[60] , \Z\R_DATA_TEMPR6[20] , 
        \Z\R_DATA_TEMPR6[21] , \Z\R_DATA_TEMPR6[38] , 
        \Z\R_DATA_TEMPR6[14] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0_DB_DETECT, 
        \Z\ACCESS_BUSY[6][0] , OR4_353_Y, \Z\R_DATA_TEMPR31[7] , 
        OR4_179_Y, OR4_33_Y, OR4_383_Y, \Z\R_DATA_TEMPR13[24] , 
        OR4_559_Y, \Z\R_DATA_TEMPR13[0] , \Z\R_DATA_TEMPR10[46] , 
        OR4_367_Y, OR4_543_Y, \Z\R_DATA_TEMPR2[44] , OR4_622_Y, 
        OR4_544_Y, OR4_48_Y, \Z\R_DATA_TEMPR21[70] , 
        \Z\R_DATA_TEMPR22[43] , \Z\R_DATA_TEMPR10[44] , 
        \Z\R_DATA_TEMPR2[42] , \Z\R_DATA_TEMPR7[66] , OR4_354_Y, 
        \Z\R_DATA_TEMPR31[38] , OR4_437_Y, \Z\R_DATA_TEMPR31[25] , 
        \Z\R_DATA_TEMPR31[27] , \Z\R_DATA_TEMPR31[30] , 
        \Z\R_DATA_TEMPR31[1] , \Z\R_DATA_TEMPR31[6] , 
        \Z\R_DATA_TEMPR31[8] , \Z\R_DATA_TEMPR31[11] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0_DB_DETECT, 
        \Z\ACCESS_BUSY[31][0] , OR4_409_Y, \Z\R_DATA_TEMPR10[68] , 
        OR4_665_Y, \Z\R_DATA_TEMPR10[62] , \Z\R_DATA_TEMPR10[74] , 
        \Z\R_DATA_TEMPR10[40] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C1_DB_DETECT, 
        \Z\ACCESS_BUSY[10][1] , OR4_177_Y, \Z\R_DATA_TEMPR2[49] , 
        OR2_22_Y, \Z\R_DATA_TEMPR21[41] , \Z\R_DATA_TEMPR7[67] , 
        \Z\R_DATA_TEMPR13[2] , \Z\R_DATA_TEMPR21[45] , 
        \Z\R_DATA_TEMPR2[53] , \Z\R_DATA_TEMPR13[33] , 
        \Z\R_DATA_TEMPR13[14] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0_DB_DETECT, 
        \Z\ACCESS_BUSY[13][0] , OR4_293_Y, \Z\R_DATA_TEMPR22[49] , 
        \Z\R_DATA_TEMPR22[41] , \Z\R_DATA_TEMPR22[73] , 
        \Z\R_DATA_TEMPR21[61] , \Z\R_DATA_TEMPR21[62] , 
        \Z\R_DATA_TEMPR21[68] , \Z\R_DATA_TEMPR21[76] , 
        \Z\R_DATA_TEMPR21[79] , \Z\R_DATA_TEMPR21[44] , 
        \Z\R_DATA_TEMPR21[51] , \Z\R_DATA_TEMPR21[53] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C1_DB_DETECT, 
        \Z\ACCESS_BUSY[21][1] , OR2_43_Y, \Z\R_DATA_TEMPR22[76] , 
        \Z\R_DATA_TEMPR7[69] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C1_DB_DETECT, 
        \Z\ACCESS_BUSY[7][1] , \Z\R_DATA_TEMPR2[74] , OR4_135_Y, 
        OR2_61_Y, \Z\R_DATA_TEMPR22[64] , \Z\R_DATA_TEMPR22[68] , 
        \Z\R_DATA_TEMPR22[74] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C1_DB_DETECT, 
        \Z\ACCESS_BUSY[22][1] , \Z\R_DATA_TEMPR2[54] , 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C1_SB_CORRECT, 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C1_DB_DETECT, 
        \Z\ACCESS_BUSY[2][1] ;
    
    OR4 OR4_700 (.A(OR4_229_Y), .B(OR4_342_Y), .C(OR4_337_Y), .D(
        OR4_455_Y), .Y(OR4_700_Y));
    OR4 OR4_399 (.A(\Z\R_DATA_TEMPR8[9] ), .B(\Z\R_DATA_TEMPR9[9] ), 
        .C(\Z\R_DATA_TEMPR10[9] ), .D(\Z\R_DATA_TEMPR11[9] ), .Y(
        OR4_399_Y));
    OR4 OR4_420 (.A(\Z\R_DATA_TEMPR28[63] ), .B(\Z\R_DATA_TEMPR29[63] )
        , .C(\Z\R_DATA_TEMPR30[63] ), .D(\Z\R_DATA_TEMPR31[63] ), .Y(
        OR4_420_Y));
    OR4 OR4_402 (.A(OR4_602_Y), .B(OR2_0_Y), .C(\Z\R_DATA_TEMPR22[74] )
        , .D(\Z\R_DATA_TEMPR23[74] ), .Y(OR4_402_Y));
    OR4 OR4_384 (.A(\Z\R_DATA_TEMPR28[1] ), .B(\Z\R_DATA_TEMPR29[1] ), 
        .C(\Z\R_DATA_TEMPR30[1] ), .D(\Z\R_DATA_TEMPR31[1] ), .Y(
        OR4_384_Y));
    OR4 OR4_373 (.A(OR4_293_Y), .B(OR2_21_Y), .C(\Z\R_DATA_TEMPR22[3] )
        , .D(\Z\R_DATA_TEMPR23[3] ), .Y(OR4_373_Y));
    OR4 \OR4_R_DATA[59]  (.A(OR4_497_Y), .B(OR4_336_Y), .C(OR4_290_Y), 
        .D(OR4_163_Y), .Y(R_DATA_c[59]));
    OR4 OR4_253 (.A(\Z\R_DATA_TEMPR24[69] ), .B(\Z\R_DATA_TEMPR25[69] )
        , .C(\Z\R_DATA_TEMPR26[69] ), .D(\Z\R_DATA_TEMPR27[69] ), .Y(
        OR4_253_Y));
    OR4 OR4_409 (.A(\Z\R_DATA_TEMPR12[33] ), .B(\Z\R_DATA_TEMPR13[33] )
        , .C(\Z\R_DATA_TEMPR14[33] ), .D(\Z\R_DATA_TEMPR15[33] ), .Y(
        OR4_409_Y));
    OR4 OR4_472 (.A(\Z\R_DATA_TEMPR24[25] ), .B(\Z\R_DATA_TEMPR25[25] )
        , .C(\Z\R_DATA_TEMPR26[25] ), .D(\Z\R_DATA_TEMPR27[25] ), .Y(
        OR4_472_Y));
    OR4 OR4_181 (.A(OR4_456_Y), .B(OR4_155_Y), .C(OR4_196_Y), .D(
        OR4_557_Y), .Y(OR4_181_Y));
    OR4 OR4_106 (.A(\Z\R_DATA_TEMPR0[54] ), .B(\Z\R_DATA_TEMPR1[54] ), 
        .C(\Z\R_DATA_TEMPR2[54] ), .D(\Z\R_DATA_TEMPR3[54] ), .Y(
        OR4_106_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[2]  (.A(CFG2_7_Y), .B(
        W_ADDR_c[13]), .C(W_EN_c), .Y(\Z\BLKX2[2] ));
    OR4 OR4_83 (.A(OR4_424_Y), .B(OR2_61_Y), .C(\Z\R_DATA_TEMPR22[68] )
        , .D(\Z\R_DATA_TEMPR23[68] ), .Y(OR4_83_Y));
    OR4 OR4_479 (.A(\Z\R_DATA_TEMPR16[8] ), .B(\Z\R_DATA_TEMPR17[8] ), 
        .C(\Z\R_DATA_TEMPR18[8] ), .D(\Z\R_DATA_TEMPR19[8] ), .Y(
        OR4_479_Y));
    OR4 OR4_138 (.A(\Z\R_DATA_TEMPR16[10] ), .B(\Z\R_DATA_TEMPR17[10] )
        , .C(\Z\R_DATA_TEMPR18[10] ), .D(\Z\R_DATA_TEMPR19[10] ), .Y(
        OR4_138_Y));
    OR4 OR4_176 (.A(OR4_340_Y), .B(OR2_74_Y), .C(
        \Z\R_DATA_TEMPR22[36] ), .D(\Z\R_DATA_TEMPR23[36] ), .Y(
        OR4_176_Y));
    OR4 OR4_610 (.A(\Z\R_DATA_TEMPR12[14] ), .B(\Z\R_DATA_TEMPR13[14] )
        , .C(\Z\R_DATA_TEMPR14[14] ), .D(\Z\R_DATA_TEMPR15[14] ), .Y(
        OR4_610_Y));
    OR2 OR2_43 (.A(\Z\R_DATA_TEMPR20[76] ), .B(\Z\R_DATA_TEMPR21[76] ), 
        .Y(OR2_43_Y));
    OR4 OR4_481 (.A(\Z\R_DATA_TEMPR28[11] ), .B(\Z\R_DATA_TEMPR29[11] )
        , .C(\Z\R_DATA_TEMPR30[11] ), .D(\Z\R_DATA_TEMPR31[11] ), .Y(
        OR4_481_Y));
    OR4 OR4_488 (.A(\Z\R_DATA_TEMPR4[38] ), .B(\Z\R_DATA_TEMPR5[38] ), 
        .C(\Z\R_DATA_TEMPR6[38] ), .D(\Z\R_DATA_TEMPR7[38] ), .Y(
        OR4_488_Y));
    OR4 OR4_308 (.A(\Z\R_DATA_TEMPR4[21] ), .B(\Z\R_DATA_TEMPR5[21] ), 
        .C(\Z\R_DATA_TEMPR6[21] ), .D(\Z\R_DATA_TEMPR7[21] ), .Y(
        OR4_308_Y));
    OR4 OR4_317 (.A(\Z\R_DATA_TEMPR4[20] ), .B(\Z\R_DATA_TEMPR5[20] ), 
        .C(\Z\R_DATA_TEMPR6[20] ), .D(\Z\R_DATA_TEMPR7[20] ), .Y(
        OR4_317_Y));
    OR4 OR4_110 (.A(\Z\R_DATA_TEMPR16[21] ), .B(\Z\R_DATA_TEMPR17[21] )
        , .C(\Z\R_DATA_TEMPR18[21] ), .D(\Z\R_DATA_TEMPR19[21] ), .Y(
        OR4_110_Y));
    OR4 OR4_658 (.A(OR4_184_Y), .B(OR4_31_Y), .C(OR4_21_Y), .D(
        OR4_460_Y), .Y(OR4_658_Y));
    OR4 OR4_378 (.A(OR4_623_Y), .B(OR4_23_Y), .C(OR4_22_Y), .D(
        OR4_135_Y), .Y(OR4_378_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%2%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C1 (
        .A_DOUT({\Z\R_DATA_TEMPR2[79] , \Z\R_DATA_TEMPR2[78] , 
        \Z\R_DATA_TEMPR2[77] , \Z\R_DATA_TEMPR2[76] , 
        \Z\R_DATA_TEMPR2[75] , \Z\R_DATA_TEMPR2[74] , 
        \Z\R_DATA_TEMPR2[73] , \Z\R_DATA_TEMPR2[72] , 
        \Z\R_DATA_TEMPR2[71] , \Z\R_DATA_TEMPR2[70] , 
        \Z\R_DATA_TEMPR2[69] , \Z\R_DATA_TEMPR2[68] , 
        \Z\R_DATA_TEMPR2[67] , \Z\R_DATA_TEMPR2[66] , 
        \Z\R_DATA_TEMPR2[65] , \Z\R_DATA_TEMPR2[64] , 
        \Z\R_DATA_TEMPR2[63] , \Z\R_DATA_TEMPR2[62] , 
        \Z\R_DATA_TEMPR2[61] , \Z\R_DATA_TEMPR2[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR2[59] , \Z\R_DATA_TEMPR2[58] , 
        \Z\R_DATA_TEMPR2[57] , \Z\R_DATA_TEMPR2[56] , 
        \Z\R_DATA_TEMPR2[55] , \Z\R_DATA_TEMPR2[54] , 
        \Z\R_DATA_TEMPR2[53] , \Z\R_DATA_TEMPR2[52] , 
        \Z\R_DATA_TEMPR2[51] , \Z\R_DATA_TEMPR2[50] , 
        \Z\R_DATA_TEMPR2[49] , \Z\R_DATA_TEMPR2[48] , 
        \Z\R_DATA_TEMPR2[47] , \Z\R_DATA_TEMPR2[46] , 
        \Z\R_DATA_TEMPR2[45] , \Z\R_DATA_TEMPR2[44] , 
        \Z\R_DATA_TEMPR2[43] , \Z\R_DATA_TEMPR2[42] , 
        \Z\R_DATA_TEMPR2[41] , \Z\R_DATA_TEMPR2[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[2][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[0] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[0] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_2 (.A(OR4_262_Y), .B(OR4_368_Y), .C(OR4_367_Y), .D(
        OR4_491_Y), .Y(OR4_2_Y));
    OR4 OR4_718 (.A(\Z\R_DATA_TEMPR4[14] ), .B(\Z\R_DATA_TEMPR5[14] ), 
        .C(\Z\R_DATA_TEMPR6[14] ), .D(\Z\R_DATA_TEMPR7[14] ), .Y(
        OR4_718_Y));
    OR2 OR2_75 (.A(\Z\R_DATA_TEMPR20[53] ), .B(\Z\R_DATA_TEMPR21[53] ), 
        .Y(OR2_75_Y));
    OR4 OR4_329 (.A(\Z\R_DATA_TEMPR24[47] ), .B(\Z\R_DATA_TEMPR25[47] )
        , .C(\Z\R_DATA_TEMPR26[47] ), .D(\Z\R_DATA_TEMPR27[47] ), .Y(
        OR4_329_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%22%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C1 (
        .A_DOUT({\Z\R_DATA_TEMPR22[79] , \Z\R_DATA_TEMPR22[78] , 
        \Z\R_DATA_TEMPR22[77] , \Z\R_DATA_TEMPR22[76] , 
        \Z\R_DATA_TEMPR22[75] , \Z\R_DATA_TEMPR22[74] , 
        \Z\R_DATA_TEMPR22[73] , \Z\R_DATA_TEMPR22[72] , 
        \Z\R_DATA_TEMPR22[71] , \Z\R_DATA_TEMPR22[70] , 
        \Z\R_DATA_TEMPR22[69] , \Z\R_DATA_TEMPR22[68] , 
        \Z\R_DATA_TEMPR22[67] , \Z\R_DATA_TEMPR22[66] , 
        \Z\R_DATA_TEMPR22[65] , \Z\R_DATA_TEMPR22[64] , 
        \Z\R_DATA_TEMPR22[63] , \Z\R_DATA_TEMPR22[62] , 
        \Z\R_DATA_TEMPR22[61] , \Z\R_DATA_TEMPR22[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR22[59] , \Z\R_DATA_TEMPR22[58] , 
        \Z\R_DATA_TEMPR22[57] , \Z\R_DATA_TEMPR22[56] , 
        \Z\R_DATA_TEMPR22[55] , \Z\R_DATA_TEMPR22[54] , 
        \Z\R_DATA_TEMPR22[53] , \Z\R_DATA_TEMPR22[52] , 
        \Z\R_DATA_TEMPR22[51] , \Z\R_DATA_TEMPR22[50] , 
        \Z\R_DATA_TEMPR22[49] , \Z\R_DATA_TEMPR22[48] , 
        \Z\R_DATA_TEMPR22[47] , \Z\R_DATA_TEMPR22[46] , 
        \Z\R_DATA_TEMPR22[45] , \Z\R_DATA_TEMPR22[44] , 
        \Z\R_DATA_TEMPR22[43] , \Z\R_DATA_TEMPR22[42] , 
        \Z\R_DATA_TEMPR22[41] , \Z\R_DATA_TEMPR22[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[22][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[5] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[5] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[29]  (.A(OR4_171_Y), .B(OR4_9_Y), .C(OR4_681_Y), 
        .D(OR4_561_Y), .Y(R_DATA_c[29]));
    OR2 OR2_63 (.A(\Z\R_DATA_TEMPR20[61] ), .B(\Z\R_DATA_TEMPR21[61] ), 
        .Y(OR2_63_Y));
    OR4 OR4_667 (.A(\Z\R_DATA_TEMPR16[75] ), .B(\Z\R_DATA_TEMPR17[75] )
        , .C(\Z\R_DATA_TEMPR18[75] ), .D(\Z\R_DATA_TEMPR19[75] ), .Y(
        OR4_667_Y));
    OR4 OR4_652 (.A(OR4_112_Y), .B(OR2_60_Y), .C(
        \Z\R_DATA_TEMPR22[64] ), .D(\Z\R_DATA_TEMPR23[64] ), .Y(
        OR4_652_Y));
    OR4 OR4_593 (.A(OR4_539_Y), .B(OR4_382_Y), .C(OR4_543_Y), .D(
        OR4_145_Y), .Y(OR4_593_Y));
    OR4 OR4_48 (.A(\Z\R_DATA_TEMPR8[74] ), .B(\Z\R_DATA_TEMPR9[74] ), 
        .C(\Z\R_DATA_TEMPR10[74] ), .D(\Z\R_DATA_TEMPR11[74] ), .Y(
        OR4_48_Y));
    OR4 OR4_589 (.A(OR4_665_Y), .B(OR4_11_Y), .C(OR4_63_Y), .D(
        OR4_16_Y), .Y(OR4_589_Y));
    OR4 OR4_109 (.A(\Z\R_DATA_TEMPR12[70] ), .B(\Z\R_DATA_TEMPR13[70] )
        , .C(\Z\R_DATA_TEMPR14[70] ), .D(\Z\R_DATA_TEMPR15[70] ), .Y(
        OR4_109_Y));
    OR2 OR2_33 (.A(\Z\R_DATA_TEMPR20[79] ), .B(\Z\R_DATA_TEMPR21[79] ), 
        .Y(OR2_33_Y));
    OR4 OR4_241 (.A(\Z\R_DATA_TEMPR24[57] ), .B(\Z\R_DATA_TEMPR25[57] )
        , .C(\Z\R_DATA_TEMPR26[57] ), .D(\Z\R_DATA_TEMPR27[57] ), .Y(
        OR4_241_Y));
    OR2 OR2_15 (.A(\Z\R_DATA_TEMPR20[44] ), .B(\Z\R_DATA_TEMPR21[44] ), 
        .Y(OR2_15_Y));
    OR4 OR4_580 (.A(\Z\R_DATA_TEMPR28[68] ), .B(\Z\R_DATA_TEMPR29[68] )
        , .C(\Z\R_DATA_TEMPR30[68] ), .D(\Z\R_DATA_TEMPR31[68] ), .Y(
        OR4_580_Y));
    OR4 OR4_81 (.A(OR4_30_Y), .B(OR4_600_Y), .C(OR4_36_Y), .D(
        OR4_364_Y), .Y(OR4_81_Y));
    OR4 OR4_118 (.A(\Z\R_DATA_TEMPR28[6] ), .B(\Z\R_DATA_TEMPR29[6] ), 
        .C(\Z\R_DATA_TEMPR30[6] ), .D(\Z\R_DATA_TEMPR31[6] ), .Y(
        OR4_118_Y));
    OR4 \OR4_R_DATA[7]  (.A(OR4_422_Y), .B(OR4_661_Y), .C(OR4_459_Y), 
        .D(OR4_353_Y), .Y(R_DATA_c[7]));
    OR4 OR4_179 (.A(\Z\R_DATA_TEMPR8[6] ), .B(\Z\R_DATA_TEMPR9[6] ), 
        .C(\Z\R_DATA_TEMPR10[6] ), .D(\Z\R_DATA_TEMPR11[6] ), .Y(
        OR4_179_Y));
    OR2 OR2_41 (.A(\Z\R_DATA_TEMPR20[62] ), .B(\Z\R_DATA_TEMPR21[62] ), 
        .Y(OR2_41_Y));
    OR4 OR4_542 (.A(\Z\R_DATA_TEMPR28[8] ), .B(\Z\R_DATA_TEMPR29[8] ), 
        .C(\Z\R_DATA_TEMPR30[8] ), .D(\Z\R_DATA_TEMPR31[8] ), .Y(
        OR4_542_Y));
    OR2 OR2_61 (.A(\Z\R_DATA_TEMPR20[68] ), .B(\Z\R_DATA_TEMPR21[68] ), 
        .Y(OR2_61_Y));
    OR4 \OR4_R_DATA[4]  (.A(OR4_556_Y), .B(OR4_136_Y), .C(OR4_246_Y), 
        .D(OR4_312_Y), .Y(R_DATA_c[4]));
    OR4 OR4_135 (.A(\Z\R_DATA_TEMPR12[41] ), .B(\Z\R_DATA_TEMPR13[41] )
        , .C(\Z\R_DATA_TEMPR14[41] ), .D(\Z\R_DATA_TEMPR15[41] ), .Y(
        OR4_135_Y));
    OR4 OR4_383 (.A(OR4_622_Y), .B(OR4_477_Y), .C(OR4_466_Y), .D(
        OR4_197_Y), .Y(OR4_383_Y));
    OR4 OR4_544 (.A(\Z\R_DATA_TEMPR0[74] ), .B(\Z\R_DATA_TEMPR1[74] ), 
        .C(\Z\R_DATA_TEMPR2[74] ), .D(\Z\R_DATA_TEMPR3[74] ), .Y(
        OR4_544_Y));
    OR4 OR4_267 (.A(\Z\R_DATA_TEMPR4[69] ), .B(\Z\R_DATA_TEMPR5[69] ), 
        .C(\Z\R_DATA_TEMPR6[69] ), .D(\Z\R_DATA_TEMPR7[69] ), .Y(
        OR4_267_Y));
    OR2 OR2_31 (.A(\Z\R_DATA_TEMPR20[51] ), .B(\Z\R_DATA_TEMPR21[51] ), 
        .Y(OR2_31_Y));
    OR4 OR4_523 (.A(\Z\R_DATA_TEMPR12[40] ), .B(\Z\R_DATA_TEMPR13[40] )
        , .C(\Z\R_DATA_TEMPR14[40] ), .D(\Z\R_DATA_TEMPR15[40] ), .Y(
        OR4_523_Y));
    OR4 OR4_437 (.A(OR4_128_Y), .B(OR2_35_Y), .C(
        \Z\R_DATA_TEMPR22[22] ), .D(\Z\R_DATA_TEMPR23[22] ), .Y(
        OR4_437_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%7%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C1 (
        .A_DOUT({\Z\R_DATA_TEMPR7[79] , \Z\R_DATA_TEMPR7[78] , 
        \Z\R_DATA_TEMPR7[77] , \Z\R_DATA_TEMPR7[76] , 
        \Z\R_DATA_TEMPR7[75] , \Z\R_DATA_TEMPR7[74] , 
        \Z\R_DATA_TEMPR7[73] , \Z\R_DATA_TEMPR7[72] , 
        \Z\R_DATA_TEMPR7[71] , \Z\R_DATA_TEMPR7[70] , 
        \Z\R_DATA_TEMPR7[69] , \Z\R_DATA_TEMPR7[68] , 
        \Z\R_DATA_TEMPR7[67] , \Z\R_DATA_TEMPR7[66] , 
        \Z\R_DATA_TEMPR7[65] , \Z\R_DATA_TEMPR7[64] , 
        \Z\R_DATA_TEMPR7[63] , \Z\R_DATA_TEMPR7[62] , 
        \Z\R_DATA_TEMPR7[61] , \Z\R_DATA_TEMPR7[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR7[59] , \Z\R_DATA_TEMPR7[58] , 
        \Z\R_DATA_TEMPR7[57] , \Z\R_DATA_TEMPR7[56] , 
        \Z\R_DATA_TEMPR7[55] , \Z\R_DATA_TEMPR7[54] , 
        \Z\R_DATA_TEMPR7[53] , \Z\R_DATA_TEMPR7[52] , 
        \Z\R_DATA_TEMPR7[51] , \Z\R_DATA_TEMPR7[50] , 
        \Z\R_DATA_TEMPR7[49] , \Z\R_DATA_TEMPR7[48] , 
        \Z\R_DATA_TEMPR7[47] , \Z\R_DATA_TEMPR7[46] , 
        \Z\R_DATA_TEMPR7[45] , \Z\R_DATA_TEMPR7[44] , 
        \Z\R_DATA_TEMPR7[43] , \Z\R_DATA_TEMPR7[42] , 
        \Z\R_DATA_TEMPR7[41] , \Z\R_DATA_TEMPR7[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[7][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[1] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[1] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_482 (.A(\Z\R_DATA_TEMPR24[68] ), .B(\Z\R_DATA_TEMPR25[68] )
        , .C(\Z\R_DATA_TEMPR26[68] ), .D(\Z\R_DATA_TEMPR27[68] ), .Y(
        OR4_482_Y));
    OR4 OR4_167 (.A(\Z\R_DATA_TEMPR8[17] ), .B(\Z\R_DATA_TEMPR9[17] ), 
        .C(\Z\R_DATA_TEMPR10[17] ), .D(\Z\R_DATA_TEMPR11[17] ), .Y(
        OR4_167_Y));
    OR4 OR4_705 (.A(OR4_146_Y), .B(OR2_43_Y), .C(
        \Z\R_DATA_TEMPR22[76] ), .D(\Z\R_DATA_TEMPR23[76] ), .Y(
        OR4_705_Y));
    OR4 OR4_607 (.A(OR4_177_Y), .B(OR4_410_Y), .C(OR4_719_Y), .D(
        OR4_296_Y), .Y(OR4_607_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%21%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C1 (
        .A_DOUT({\Z\R_DATA_TEMPR21[79] , \Z\R_DATA_TEMPR21[78] , 
        \Z\R_DATA_TEMPR21[77] , \Z\R_DATA_TEMPR21[76] , 
        \Z\R_DATA_TEMPR21[75] , \Z\R_DATA_TEMPR21[74] , 
        \Z\R_DATA_TEMPR21[73] , \Z\R_DATA_TEMPR21[72] , 
        \Z\R_DATA_TEMPR21[71] , \Z\R_DATA_TEMPR21[70] , 
        \Z\R_DATA_TEMPR21[69] , \Z\R_DATA_TEMPR21[68] , 
        \Z\R_DATA_TEMPR21[67] , \Z\R_DATA_TEMPR21[66] , 
        \Z\R_DATA_TEMPR21[65] , \Z\R_DATA_TEMPR21[64] , 
        \Z\R_DATA_TEMPR21[63] , \Z\R_DATA_TEMPR21[62] , 
        \Z\R_DATA_TEMPR21[61] , \Z\R_DATA_TEMPR21[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR21[59] , \Z\R_DATA_TEMPR21[58] , 
        \Z\R_DATA_TEMPR21[57] , \Z\R_DATA_TEMPR21[56] , 
        \Z\R_DATA_TEMPR21[55] , \Z\R_DATA_TEMPR21[54] , 
        \Z\R_DATA_TEMPR21[53] , \Z\R_DATA_TEMPR21[52] , 
        \Z\R_DATA_TEMPR21[51] , \Z\R_DATA_TEMPR21[50] , 
        \Z\R_DATA_TEMPR21[49] , \Z\R_DATA_TEMPR21[48] , 
        \Z\R_DATA_TEMPR21[47] , \Z\R_DATA_TEMPR21[46] , 
        \Z\R_DATA_TEMPR21[45] , \Z\R_DATA_TEMPR21[44] , 
        \Z\R_DATA_TEMPR21[43] , \Z\R_DATA_TEMPR21[42] , 
        \Z\R_DATA_TEMPR21[41] , \Z\R_DATA_TEMPR21[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[21][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[5] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[5] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_489 (.A(\Z\R_DATA_TEMPR12[77] ), .B(\Z\R_DATA_TEMPR13[77] )
        , .C(\Z\R_DATA_TEMPR14[77] ), .D(\Z\R_DATA_TEMPR15[77] ), .Y(
        OR4_489_Y));
    OR4 OR4_706 (.A(\Z\R_DATA_TEMPR24[11] ), .B(\Z\R_DATA_TEMPR25[11] )
        , .C(\Z\R_DATA_TEMPR26[11] ), .D(\Z\R_DATA_TEMPR27[11] ), .Y(
        OR4_706_Y));
    OR4 OR4_186 (.A(\Z\R_DATA_TEMPR24[67] ), .B(\Z\R_DATA_TEMPR25[67] )
        , .C(\Z\R_DATA_TEMPR26[67] ), .D(\Z\R_DATA_TEMPR27[67] ), .Y(
        OR4_186_Y));
    OR4 OR4_677 (.A(OR4_427_Y), .B(OR2_68_Y), .C(\Z\R_DATA_TEMPR22[1] )
        , .D(\Z\R_DATA_TEMPR23[1] ), .Y(OR4_677_Y));
    OR4 OR4_341 (.A(OR4_559_Y), .B(OR2_22_Y), .C(
        \Z\R_DATA_TEMPR22[41] ), .D(\Z\R_DATA_TEMPR23[41] ), .Y(
        OR4_341_Y));
    OR4 OR4_235 (.A(OR4_89_Y), .B(OR2_57_Y), .C(\Z\R_DATA_TEMPR22[73] )
        , .D(\Z\R_DATA_TEMPR23[73] ), .Y(OR4_235_Y));
    OR2 OR2_29 (.A(\Z\R_DATA_TEMPR20[18] ), .B(\Z\R_DATA_TEMPR21[18] ), 
        .Y(OR2_29_Y));
    OR4 OR4_264 (.A(\Z\R_DATA_TEMPR28[30] ), .B(\Z\R_DATA_TEMPR29[30] )
        , .C(\Z\R_DATA_TEMPR30[30] ), .D(\Z\R_DATA_TEMPR31[30] ), .Y(
        OR4_264_Y));
    OR4 OR4_656 (.A(\Z\R_DATA_TEMPR0[12] ), .B(\Z\R_DATA_TEMPR1[12] ), 
        .C(\Z\R_DATA_TEMPR2[12] ), .D(\Z\R_DATA_TEMPR3[12] ), .Y(
        OR4_656_Y));
    OR4 OR4_440 (.A(OR4_41_Y), .B(OR2_48_Y), .C(\Z\R_DATA_TEMPR22[49] )
        , .D(\Z\R_DATA_TEMPR23[49] ), .Y(OR4_440_Y));
    OR4 OR4_293 (.A(\Z\R_DATA_TEMPR16[3] ), .B(\Z\R_DATA_TEMPR17[3] ), 
        .C(\Z\R_DATA_TEMPR18[3] ), .D(\Z\R_DATA_TEMPR19[3] ), .Y(
        OR4_293_Y));
    OR4 OR4_388 (.A(\Z\R_DATA_TEMPR28[66] ), .B(\Z\R_DATA_TEMPR29[66] )
        , .C(\Z\R_DATA_TEMPR30[66] ), .D(\Z\R_DATA_TEMPR31[66] ), .Y(
        OR4_388_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%13%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0 (
        .A_DOUT({\Z\R_DATA_TEMPR13[39] , \Z\R_DATA_TEMPR13[38] , 
        \Z\R_DATA_TEMPR13[37] , \Z\R_DATA_TEMPR13[36] , 
        \Z\R_DATA_TEMPR13[35] , \Z\R_DATA_TEMPR13[34] , 
        \Z\R_DATA_TEMPR13[33] , \Z\R_DATA_TEMPR13[32] , 
        \Z\R_DATA_TEMPR13[31] , \Z\R_DATA_TEMPR13[30] , 
        \Z\R_DATA_TEMPR13[29] , \Z\R_DATA_TEMPR13[28] , 
        \Z\R_DATA_TEMPR13[27] , \Z\R_DATA_TEMPR13[26] , 
        \Z\R_DATA_TEMPR13[25] , \Z\R_DATA_TEMPR13[24] , 
        \Z\R_DATA_TEMPR13[23] , \Z\R_DATA_TEMPR13[22] , 
        \Z\R_DATA_TEMPR13[21] , \Z\R_DATA_TEMPR13[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR13[19] , \Z\R_DATA_TEMPR13[18] , 
        \Z\R_DATA_TEMPR13[17] , \Z\R_DATA_TEMPR13[16] , 
        \Z\R_DATA_TEMPR13[15] , \Z\R_DATA_TEMPR13[14] , 
        \Z\R_DATA_TEMPR13[13] , \Z\R_DATA_TEMPR13[12] , 
        \Z\R_DATA_TEMPR13[11] , \Z\R_DATA_TEMPR13[10] , 
        \Z\R_DATA_TEMPR13[9] , \Z\R_DATA_TEMPR13[8] , 
        \Z\R_DATA_TEMPR13[7] , \Z\R_DATA_TEMPR13[6] , 
        \Z\R_DATA_TEMPR13[5] , \Z\R_DATA_TEMPR13[4] , 
        \Z\R_DATA_TEMPR13[3] , \Z\R_DATA_TEMPR13[2] , 
        \Z\R_DATA_TEMPR13[1] , \Z\R_DATA_TEMPR13[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[13][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[3] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[3] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_115 (.A(OR4_404_Y), .B(OR4_94_Y), .C(OR4_127_Y), .D(
        OR4_503_Y), .Y(OR4_115_Y));
    OR4 OR4_66 (.A(OR4_386_Y), .B(OR2_55_Y), .C(\Z\R_DATA_TEMPR22[19] )
        , .D(\Z\R_DATA_TEMPR23[19] ), .Y(OR4_66_Y));
    OR4 OR4_433 (.A(OR4_331_Y), .B(OR2_71_Y), .C(
        \Z\R_DATA_TEMPR22[27] ), .D(\Z\R_DATA_TEMPR23[27] ), .Y(
        OR4_433_Y));
    OR4 OR4_417 (.A(\Z\R_DATA_TEMPR24[9] ), .B(\Z\R_DATA_TEMPR25[9] ), 
        .C(\Z\R_DATA_TEMPR26[9] ), .D(\Z\R_DATA_TEMPR27[9] ), .Y(
        OR4_417_Y));
    OR4 OR4_631 (.A(\Z\R_DATA_TEMPR16[14] ), .B(\Z\R_DATA_TEMPR17[14] )
        , .C(\Z\R_DATA_TEMPR18[14] ), .D(\Z\R_DATA_TEMPR19[14] ), .Y(
        OR4_631_Y));
    OR4 OR4_365 (.A(\Z\R_DATA_TEMPR8[38] ), .B(\Z\R_DATA_TEMPR9[38] ), 
        .C(\Z\R_DATA_TEMPR10[38] ), .D(\Z\R_DATA_TEMPR11[38] ), .Y(
        OR4_365_Y));
    CFG2 #( .INIT(4'h1) )  CFG2_4 (.A(W_ADDR_c[12]), .B(W_ADDR_c[11]), 
        .Y(CFG2_4_Y));
    OR4 OR4_238 (.A(\Z\R_DATA_TEMPR0[53] ), .B(\Z\R_DATA_TEMPR1[53] ), 
        .C(\Z\R_DATA_TEMPR2[53] ), .D(\Z\R_DATA_TEMPR3[53] ), .Y(
        OR4_238_Y));
    OR2 OR2_8 (.A(\Z\R_DATA_TEMPR20[45] ), .B(\Z\R_DATA_TEMPR21[45] ), 
        .Y(OR2_8_Y));
    OR4 \OR4_R_DATA[52]  (.A(OR4_62_Y), .B(OR4_44_Y), .C(OR4_671_Y), 
        .D(OR4_344_Y), .Y(R_DATA_c[52]));
    OR4 OR4_189 (.A(OR4_59_Y), .B(OR4_226_Y), .C(OR4_295_Y), .D(
        OR4_93_Y), .Y(OR4_189_Y));
    OR4 OR4_0 (.A(\Z\R_DATA_TEMPR8[62] ), .B(\Z\R_DATA_TEMPR9[62] ), 
        .C(\Z\R_DATA_TEMPR10[62] ), .D(\Z\R_DATA_TEMPR11[62] ), .Y(
        OR4_0_Y));
    OR4 OR4_207 (.A(\Z\R_DATA_TEMPR8[40] ), .B(\Z\R_DATA_TEMPR9[40] ), 
        .C(\Z\R_DATA_TEMPR10[40] ), .D(\Z\R_DATA_TEMPR11[40] ), .Y(
        OR4_207_Y));
    OR4 OR4_215 (.A(\Z\R_DATA_TEMPR12[2] ), .B(\Z\R_DATA_TEMPR13[2] ), 
        .C(\Z\R_DATA_TEMPR14[2] ), .D(\Z\R_DATA_TEMPR15[2] ), .Y(
        OR4_215_Y));
    OR4 OR4_107 (.A(OR4_321_Y), .B(OR4_575_Y), .C(OR4_516_Y), .D(
        OR4_228_Y), .Y(OR4_107_Y));
    OR4 OR4_277 (.A(OR4_517_Y), .B(OR4_643_Y), .C(OR4_640_Y), .D(
        OR4_33_Y), .Y(OR4_277_Y));
    OR4 OR4_95 (.A(\Z\R_DATA_TEMPR4[67] ), .B(\Z\R_DATA_TEMPR5[67] ), 
        .C(\Z\R_DATA_TEMPR6[67] ), .D(\Z\R_DATA_TEMPR7[67] ), .Y(
        OR4_95_Y));
    OR4 OR4_698 (.A(OR4_74_Y), .B(OR2_40_Y), .C(\Z\R_DATA_TEMPR22[20] )
        , .D(\Z\R_DATA_TEMPR23[20] ), .Y(OR4_698_Y));
    OR2 OR2_22 (.A(\Z\R_DATA_TEMPR20[41] ), .B(\Z\R_DATA_TEMPR21[41] ), 
        .Y(OR2_22_Y));
    OR4 OR4_177 (.A(\Z\R_DATA_TEMPR0[49] ), .B(\Z\R_DATA_TEMPR1[49] ), 
        .C(\Z\R_DATA_TEMPR2[49] ), .D(\Z\R_DATA_TEMPR3[49] ), .Y(
        OR4_177_Y));
    OR2 OR2_79 (.A(\Z\R_DATA_TEMPR20[29] ), .B(\Z\R_DATA_TEMPR21[29] ), 
        .Y(OR2_79_Y));
    OR4 \OR4_R_DATA[34]  (.A(OR4_122_Y), .B(OR4_604_Y), .C(OR4_243_Y), 
        .D(OR4_547_Y), .Y(R_DATA_c[34]));
    OR4 OR4_349 (.A(\Z\R_DATA_TEMPR28[50] ), .B(\Z\R_DATA_TEMPR29[50] )
        , .C(\Z\R_DATA_TEMPR30[50] ), .D(\Z\R_DATA_TEMPR31[50] ), .Y(
        OR4_349_Y));
    OR4 OR4_692 (.A(\Z\R_DATA_TEMPR28[27] ), .B(\Z\R_DATA_TEMPR29[27] )
        , .C(\Z\R_DATA_TEMPR30[27] ), .D(\Z\R_DATA_TEMPR31[27] ), .Y(
        OR4_692_Y));
    OR4 OR4_703 (.A(\Z\R_DATA_TEMPR0[30] ), .B(\Z\R_DATA_TEMPR1[30] ), 
        .C(\Z\R_DATA_TEMPR2[30] ), .D(\Z\R_DATA_TEMPR3[30] ), .Y(
        OR4_703_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%10%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C1 (
        .A_DOUT({\Z\R_DATA_TEMPR10[79] , \Z\R_DATA_TEMPR10[78] , 
        \Z\R_DATA_TEMPR10[77] , \Z\R_DATA_TEMPR10[76] , 
        \Z\R_DATA_TEMPR10[75] , \Z\R_DATA_TEMPR10[74] , 
        \Z\R_DATA_TEMPR10[73] , \Z\R_DATA_TEMPR10[72] , 
        \Z\R_DATA_TEMPR10[71] , \Z\R_DATA_TEMPR10[70] , 
        \Z\R_DATA_TEMPR10[69] , \Z\R_DATA_TEMPR10[68] , 
        \Z\R_DATA_TEMPR10[67] , \Z\R_DATA_TEMPR10[66] , 
        \Z\R_DATA_TEMPR10[65] , \Z\R_DATA_TEMPR10[64] , 
        \Z\R_DATA_TEMPR10[63] , \Z\R_DATA_TEMPR10[62] , 
        \Z\R_DATA_TEMPR10[61] , \Z\R_DATA_TEMPR10[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR10[59] , \Z\R_DATA_TEMPR10[58] , 
        \Z\R_DATA_TEMPR10[57] , \Z\R_DATA_TEMPR10[56] , 
        \Z\R_DATA_TEMPR10[55] , \Z\R_DATA_TEMPR10[54] , 
        \Z\R_DATA_TEMPR10[53] , \Z\R_DATA_TEMPR10[52] , 
        \Z\R_DATA_TEMPR10[51] , \Z\R_DATA_TEMPR10[50] , 
        \Z\R_DATA_TEMPR10[49] , \Z\R_DATA_TEMPR10[48] , 
        \Z\R_DATA_TEMPR10[47] , \Z\R_DATA_TEMPR10[46] , 
        \Z\R_DATA_TEMPR10[45] , \Z\R_DATA_TEMPR10[44] , 
        \Z\R_DATA_TEMPR10[43] , \Z\R_DATA_TEMPR10[42] , 
        \Z\R_DATA_TEMPR10[41] , \Z\R_DATA_TEMPR10[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[10][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[2] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[2] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_223 (.A(\Z\R_DATA_TEMPR0[17] ), .B(\Z\R_DATA_TEMPR1[17] ), 
        .C(\Z\R_DATA_TEMPR2[17] ), .D(\Z\R_DATA_TEMPR3[17] ), .Y(
        OR4_223_Y));
    OR4 OR4_354 (.A(\Z\R_DATA_TEMPR0[35] ), .B(\Z\R_DATA_TEMPR1[35] ), 
        .C(\Z\R_DATA_TEMPR2[35] ), .D(\Z\R_DATA_TEMPR3[35] ), .Y(
        OR4_354_Y));
    OR4 OR4_204 (.A(\Z\R_DATA_TEMPR0[15] ), .B(\Z\R_DATA_TEMPR1[15] ), 
        .C(\Z\R_DATA_TEMPR2[15] ), .D(\Z\R_DATA_TEMPR3[15] ), .Y(
        OR4_204_Y));
    OR2 OR2_19 (.A(\Z\R_DATA_TEMPR20[6] ), .B(\Z\R_DATA_TEMPR21[6] ), 
        .Y(OR2_19_Y));
    OR4 OR4_665 (.A(\Z\R_DATA_TEMPR0[1] ), .B(\Z\R_DATA_TEMPR1[1] ), 
        .C(\Z\R_DATA_TEMPR2[1] ), .D(\Z\R_DATA_TEMPR3[1] ), .Y(
        OR4_665_Y));
    OR4 OR4_413 (.A(\Z\R_DATA_TEMPR8[68] ), .B(\Z\R_DATA_TEMPR9[68] ), 
        .C(\Z\R_DATA_TEMPR10[68] ), .D(\Z\R_DATA_TEMPR11[68] ), .Y(
        OR4_413_Y));
    OR4 OR4_611 (.A(OR4_116_Y), .B(OR4_709_Y), .C(OR4_693_Y), .D(
        OR4_409_Y), .Y(OR4_611_Y));
    OR4 OR4_274 (.A(\Z\R_DATA_TEMPR28[25] ), .B(\Z\R_DATA_TEMPR29[25] )
        , .C(\Z\R_DATA_TEMPR30[25] ), .D(\Z\R_DATA_TEMPR31[25] ), .Y(
        OR4_274_Y));
    OR4 OR4_151 (.A(\Z\R_DATA_TEMPR0[27] ), .B(\Z\R_DATA_TEMPR1[27] ), 
        .C(\Z\R_DATA_TEMPR2[27] ), .D(\Z\R_DATA_TEMPR3[27] ), .Y(
        OR4_151_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%31%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0 (
        .A_DOUT({\Z\R_DATA_TEMPR31[39] , \Z\R_DATA_TEMPR31[38] , 
        \Z\R_DATA_TEMPR31[37] , \Z\R_DATA_TEMPR31[36] , 
        \Z\R_DATA_TEMPR31[35] , \Z\R_DATA_TEMPR31[34] , 
        \Z\R_DATA_TEMPR31[33] , \Z\R_DATA_TEMPR31[32] , 
        \Z\R_DATA_TEMPR31[31] , \Z\R_DATA_TEMPR31[30] , 
        \Z\R_DATA_TEMPR31[29] , \Z\R_DATA_TEMPR31[28] , 
        \Z\R_DATA_TEMPR31[27] , \Z\R_DATA_TEMPR31[26] , 
        \Z\R_DATA_TEMPR31[25] , \Z\R_DATA_TEMPR31[24] , 
        \Z\R_DATA_TEMPR31[23] , \Z\R_DATA_TEMPR31[22] , 
        \Z\R_DATA_TEMPR31[21] , \Z\R_DATA_TEMPR31[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR31[19] , \Z\R_DATA_TEMPR31[18] , 
        \Z\R_DATA_TEMPR31[17] , \Z\R_DATA_TEMPR31[16] , 
        \Z\R_DATA_TEMPR31[15] , \Z\R_DATA_TEMPR31[14] , 
        \Z\R_DATA_TEMPR31[13] , \Z\R_DATA_TEMPR31[12] , 
        \Z\R_DATA_TEMPR31[11] , \Z\R_DATA_TEMPR31[10] , 
        \Z\R_DATA_TEMPR31[9] , \Z\R_DATA_TEMPR31[8] , 
        \Z\R_DATA_TEMPR31[7] , \Z\R_DATA_TEMPR31[6] , 
        \Z\R_DATA_TEMPR31[5] , \Z\R_DATA_TEMPR31[4] , 
        \Z\R_DATA_TEMPR31[3] , \Z\R_DATA_TEMPR31[2] , 
        \Z\R_DATA_TEMPR31[1] , \Z\R_DATA_TEMPR31[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[31][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[7] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[7] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_218 (.A(OR4_492_Y), .B(OR4_7_Y), .C(OR4_318_Y), .D(
        OR4_617_Y), .Y(OR4_218_Y));
    OR4 \OR4_R_DATA[22]  (.A(OR4_462_Y), .B(OR4_437_Y), .C(OR4_339_Y), 
        .D(OR4_18_Y), .Y(R_DATA_c[22]));
    OR4 \OR4_R_DATA[53]  (.A(OR4_712_Y), .B(OR4_521_Y), .C(OR4_493_Y), 
        .D(OR4_470_Y), .Y(R_DATA_c[53]));
    OR4 OR4_60 (.A(\Z\R_DATA_TEMPR24[14] ), .B(\Z\R_DATA_TEMPR25[14] ), 
        .C(\Z\R_DATA_TEMPR26[14] ), .D(\Z\R_DATA_TEMPR27[14] ), .Y(
        OR4_60_Y));
    OR4 OR4_531 (.A(\Z\R_DATA_TEMPR28[38] ), .B(\Z\R_DATA_TEMPR29[38] )
        , .C(\Z\R_DATA_TEMPR30[38] ), .D(\Z\R_DATA_TEMPR31[38] ), .Y(
        OR4_531_Y));
    OR4 OR4_67 (.A(OR4_354_Y), .B(OR4_50_Y), .C(OR4_77_Y), .D(
        OR4_449_Y), .Y(OR4_67_Y));
    OR4 OR4_687 (.A(\Z\R_DATA_TEMPR4[66] ), .B(\Z\R_DATA_TEMPR5[66] ), 
        .C(\Z\R_DATA_TEMPR6[66] ), .D(\Z\R_DATA_TEMPR7[66] ), .Y(
        OR4_687_Y));
    OR4 OR4_305 (.A(\Z\R_DATA_TEMPR0[42] ), .B(\Z\R_DATA_TEMPR1[42] ), 
        .C(\Z\R_DATA_TEMPR2[42] ), .D(\Z\R_DATA_TEMPR3[42] ), .Y(
        OR4_305_Y));
    OR4 OR4_451 (.A(\Z\R_DATA_TEMPR8[44] ), .B(\Z\R_DATA_TEMPR9[44] ), 
        .C(\Z\R_DATA_TEMPR10[44] ), .D(\Z\R_DATA_TEMPR11[44] ), .Y(
        OR4_451_Y));
    OR4 OR4_458 (.A(\Z\R_DATA_TEMPR0[29] ), .B(\Z\R_DATA_TEMPR1[29] ), 
        .C(\Z\R_DATA_TEMPR2[29] ), .D(\Z\R_DATA_TEMPR3[29] ), .Y(
        OR4_458_Y));
    OR4 OR4_628 (.A(OR4_496_Y), .B(OR2_70_Y), .C(
        \Z\R_DATA_TEMPR22[43] ), .D(\Z\R_DATA_TEMPR23[43] ), .Y(
        OR4_628_Y));
    OR4 OR4_375 (.A(\Z\R_DATA_TEMPR16[9] ), .B(\Z\R_DATA_TEMPR17[9] ), 
        .C(\Z\R_DATA_TEMPR18[9] ), .D(\Z\R_DATA_TEMPR19[9] ), .Y(
        OR4_375_Y));
    OR2 OR2_72 (.A(\Z\R_DATA_TEMPR20[70] ), .B(\Z\R_DATA_TEMPR21[70] ), 
        .Y(OR2_72_Y));
    OR4 OR4_660 (.A(OR4_544_Y), .B(OR4_699_Y), .C(OR4_48_Y), .D(
        OR4_581_Y), .Y(OR4_660_Y));
    OR4 OR4_622 (.A(\Z\R_DATA_TEMPR0[23] ), .B(\Z\R_DATA_TEMPR1[23] ), 
        .C(\Z\R_DATA_TEMPR2[23] ), .D(\Z\R_DATA_TEMPR3[23] ), .Y(
        OR4_622_Y));
    OR4 OR4_232 (.A(\Z\R_DATA_TEMPR0[44] ), .B(\Z\R_DATA_TEMPR1[44] ), 
        .C(\Z\R_DATA_TEMPR2[44] ), .D(\Z\R_DATA_TEMPR3[44] ), .Y(
        OR4_232_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[4]  (.A(CFG2_3_Y), .B(
        R_ADDR_c[13]), .C(R_EN_c), .Y(\Z\BLKY2[4] ));
    OR4 \OR4_R_DATA[15]  (.A(OR4_636_Y), .B(OR4_265_Y), .C(OR4_535_Y), 
        .D(OR4_320_Y), .Y(R_DATA_c[15]));
    OR4 OR4_543 (.A(\Z\R_DATA_TEMPR8[10] ), .B(\Z\R_DATA_TEMPR9[10] ), 
        .C(\Z\R_DATA_TEMPR10[10] ), .D(\Z\R_DATA_TEMPR11[10] ), .Y(
        OR4_543_Y));
    OR4 OR4_45 (.A(\Z\R_DATA_TEMPR28[72] ), .B(\Z\R_DATA_TEMPR29[72] ), 
        .C(\Z\R_DATA_TEMPR30[72] ), .D(\Z\R_DATA_TEMPR31[72] ), .Y(
        OR4_45_Y));
    OR4 OR4_367 (.A(\Z\R_DATA_TEMPR8[11] ), .B(\Z\R_DATA_TEMPR9[11] ), 
        .C(\Z\R_DATA_TEMPR10[11] ), .D(\Z\R_DATA_TEMPR11[11] ), .Y(
        OR4_367_Y));
    OR4 OR4_160 (.A(\Z\R_DATA_TEMPR8[46] ), .B(\Z\R_DATA_TEMPR9[46] ), 
        .C(\Z\R_DATA_TEMPR10[46] ), .D(\Z\R_DATA_TEMPR11[46] ), .Y(
        OR4_160_Y));
    OR2 OR2_12 (.A(\Z\R_DATA_TEMPR20[10] ), .B(\Z\R_DATA_TEMPR21[10] ), 
        .Y(OR2_12_Y));
    OR4 OR4_702 (.A(\Z\R_DATA_TEMPR12[0] ), .B(\Z\R_DATA_TEMPR13[0] ), 
        .C(\Z\R_DATA_TEMPR14[0] ), .D(\Z\R_DATA_TEMPR15[0] ), .Y(
        OR4_702_Y));
    OR4 OR4_559 (.A(\Z\R_DATA_TEMPR16[41] ), .B(\Z\R_DATA_TEMPR17[41] )
        , .C(\Z\R_DATA_TEMPR18[41] ), .D(\Z\R_DATA_TEMPR19[41] ), .Y(
        OR4_559_Y));
    OR4 \OR4_R_DATA[23]  (.A(OR4_383_Y), .B(OR4_206_Y), .C(OR4_164_Y), 
        .D(OR4_139_Y), .Y(R_DATA_c[23]));
    OR4 OR4_550 (.A(\Z\R_DATA_TEMPR12[24] ), .B(\Z\R_DATA_TEMPR13[24] )
        , .C(\Z\R_DATA_TEMPR14[24] ), .D(\Z\R_DATA_TEMPR15[24] ), .Y(
        OR4_550_Y));
    OR4 OR4_330 (.A(OR4_684_Y), .B(OR4_471_Y), .C(OR4_509_Y), .D(
        OR4_645_Y), .Y(OR4_330_Y));
    OR4 OR4_605 (.A(OR4_161_Y), .B(OR4_583_Y), .C(OR4_615_Y), .D(
        OR4_269_Y), .Y(OR4_605_Y));
    OR4 OR4_511 (.A(\Z\R_DATA_TEMPR0[24] ), .B(\Z\R_DATA_TEMPR1[24] ), 
        .C(\Z\R_DATA_TEMPR2[24] ), .D(\Z\R_DATA_TEMPR3[24] ), .Y(
        OR4_511_Y));
    OR4 OR4_696 (.A(\Z\R_DATA_TEMPR0[7] ), .B(\Z\R_DATA_TEMPR1[7] ), 
        .C(\Z\R_DATA_TEMPR2[7] ), .D(\Z\R_DATA_TEMPR3[7] ), .Y(
        OR4_696_Y));
    OR4 OR4_675 (.A(\Z\R_DATA_TEMPR8[32] ), .B(\Z\R_DATA_TEMPR9[32] ), 
        .C(\Z\R_DATA_TEMPR10[32] ), .D(\Z\R_DATA_TEMPR11[32] ), .Y(
        OR4_675_Y));
    OR4 OR4_86 (.A(\Z\R_DATA_TEMPR8[4] ), .B(\Z\R_DATA_TEMPR9[4] ), .C(
        \Z\R_DATA_TEMPR10[4] ), .D(\Z\R_DATA_TEMPR11[4] ), .Y(OR4_86_Y)
        );
    OR4 OR4_287 (.A(\Z\R_DATA_TEMPR12[46] ), .B(\Z\R_DATA_TEMPR13[46] )
        , .C(\Z\R_DATA_TEMPR14[46] ), .D(\Z\R_DATA_TEMPR15[46] ), .Y(
        OR4_287_Y));
    OR4 OR4_33 (.A(\Z\R_DATA_TEMPR12[51] ), .B(\Z\R_DATA_TEMPR13[51] ), 
        .C(\Z\R_DATA_TEMPR14[51] ), .D(\Z\R_DATA_TEMPR15[51] ), .Y(
        OR4_33_Y));
    OR4 OR4_168 (.A(OR4_92_Y), .B(OR4_327_Y), .C(OR4_179_Y), .D(
        OR4_174_Y), .Y(OR4_168_Y));
    OR4 OR4_187 (.A(\Z\R_DATA_TEMPR16[11] ), .B(\Z\R_DATA_TEMPR17[11] )
        , .C(\Z\R_DATA_TEMPR18[11] ), .D(\Z\R_DATA_TEMPR19[11] ), .Y(
        OR4_187_Y));
    OR2 OR2_46 (.A(\Z\R_DATA_TEMPR20[2] ), .B(\Z\R_DATA_TEMPR21[2] ), 
        .Y(OR2_46_Y));
    OR4 OR4_212 (.A(\Z\R_DATA_TEMPR8[18] ), .B(\Z\R_DATA_TEMPR9[18] ), 
        .C(\Z\R_DATA_TEMPR10[18] ), .D(\Z\R_DATA_TEMPR11[18] ), .Y(
        OR4_212_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%6%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0 (
        .A_DOUT({\Z\R_DATA_TEMPR6[39] , \Z\R_DATA_TEMPR6[38] , 
        \Z\R_DATA_TEMPR6[37] , \Z\R_DATA_TEMPR6[36] , 
        \Z\R_DATA_TEMPR6[35] , \Z\R_DATA_TEMPR6[34] , 
        \Z\R_DATA_TEMPR6[33] , \Z\R_DATA_TEMPR6[32] , 
        \Z\R_DATA_TEMPR6[31] , \Z\R_DATA_TEMPR6[30] , 
        \Z\R_DATA_TEMPR6[29] , \Z\R_DATA_TEMPR6[28] , 
        \Z\R_DATA_TEMPR6[27] , \Z\R_DATA_TEMPR6[26] , 
        \Z\R_DATA_TEMPR6[25] , \Z\R_DATA_TEMPR6[24] , 
        \Z\R_DATA_TEMPR6[23] , \Z\R_DATA_TEMPR6[22] , 
        \Z\R_DATA_TEMPR6[21] , \Z\R_DATA_TEMPR6[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR6[19] , \Z\R_DATA_TEMPR6[18] , 
        \Z\R_DATA_TEMPR6[17] , \Z\R_DATA_TEMPR6[16] , 
        \Z\R_DATA_TEMPR6[15] , \Z\R_DATA_TEMPR6[14] , 
        \Z\R_DATA_TEMPR6[13] , \Z\R_DATA_TEMPR6[12] , 
        \Z\R_DATA_TEMPR6[11] , \Z\R_DATA_TEMPR6[10] , 
        \Z\R_DATA_TEMPR6[9] , \Z\R_DATA_TEMPR6[8] , 
        \Z\R_DATA_TEMPR6[7] , \Z\R_DATA_TEMPR6[6] , 
        \Z\R_DATA_TEMPR6[5] , \Z\R_DATA_TEMPR6[4] , 
        \Z\R_DATA_TEMPR6[3] , \Z\R_DATA_TEMPR6[2] , 
        \Z\R_DATA_TEMPR6[1] , \Z\R_DATA_TEMPR6[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[6][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[1] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[1] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_353 (.A(\Z\R_DATA_TEMPR28[7] ), .B(\Z\R_DATA_TEMPR29[7] ), 
        .C(\Z\R_DATA_TEMPR30[7] ), .D(\Z\R_DATA_TEMPR31[7] ), .Y(
        OR4_353_Y));
    OR4 \OR4_R_DATA[45]  (.A(OR4_282_Y), .B(OR4_627_Y), .C(OR4_194_Y), 
        .D(OR4_707_Y), .Y(R_DATA_c[45]));
    OR4 OR4_600 (.A(\Z\R_DATA_TEMPR4[60] ), .B(\Z\R_DATA_TEMPR5[60] ), 
        .C(\Z\R_DATA_TEMPR6[60] ), .D(\Z\R_DATA_TEMPR7[60] ), .Y(
        OR4_600_Y));
    OR4 OR4_452 (.A(\Z\R_DATA_TEMPR24[0] ), .B(\Z\R_DATA_TEMPR25[0] ), 
        .C(\Z\R_DATA_TEMPR26[0] ), .D(\Z\R_DATA_TEMPR27[0] ), .Y(
        OR4_452_Y));
    OR4 OR4_310 (.A(\Z\R_DATA_TEMPR12[32] ), .B(\Z\R_DATA_TEMPR13[32] )
        , .C(\Z\R_DATA_TEMPR14[32] ), .D(\Z\R_DATA_TEMPR15[32] ), .Y(
        OR4_310_Y));
    OR4 OR4_284 (.A(\Z\R_DATA_TEMPR12[15] ), .B(\Z\R_DATA_TEMPR13[15] )
        , .C(\Z\R_DATA_TEMPR14[15] ), .D(\Z\R_DATA_TEMPR15[15] ), .Y(
        OR4_284_Y));
    OR4 OR4_5 (.A(\Z\R_DATA_TEMPR12[67] ), .B(\Z\R_DATA_TEMPR13[67] ), 
        .C(\Z\R_DATA_TEMPR14[67] ), .D(\Z\R_DATA_TEMPR15[67] ), .Y(
        OR4_5_Y));
    OR4 OR4_670 (.A(OR4_563_Y), .B(OR2_58_Y), .C(
        \Z\R_DATA_TEMPR22[37] ), .D(\Z\R_DATA_TEMPR23[37] ), .Y(
        OR4_670_Y));
    OR2 OR2_66 (.A(\Z\R_DATA_TEMPR20[56] ), .B(\Z\R_DATA_TEMPR21[56] ), 
        .Y(OR2_66_Y));
    VCC VCC_Z (.Y(VCC));
    OR4 OR4_459 (.A(\Z\R_DATA_TEMPR24[7] ), .B(\Z\R_DATA_TEMPR25[7] ), 
        .C(\Z\R_DATA_TEMPR26[7] ), .D(\Z\R_DATA_TEMPR27[7] ), .Y(
        OR4_459_Y));
    OR4 OR4_307 (.A(\Z\R_DATA_TEMPR8[21] ), .B(\Z\R_DATA_TEMPR9[21] ), 
        .C(\Z\R_DATA_TEMPR10[21] ), .D(\Z\R_DATA_TEMPR11[21] ), .Y(
        OR4_307_Y));
    OR4 OR4_100 (.A(\Z\R_DATA_TEMPR0[8] ), .B(\Z\R_DATA_TEMPR1[8] ), 
        .C(\Z\R_DATA_TEMPR2[8] ), .D(\Z\R_DATA_TEMPR3[8] ), .Y(
        OR4_100_Y));
    OR4 OR4_99 (.A(\Z\R_DATA_TEMPR16[0] ), .B(\Z\R_DATA_TEMPR17[0] ), 
        .C(\Z\R_DATA_TEMPR18[0] ), .D(\Z\R_DATA_TEMPR19[0] ), .Y(
        OR4_99_Y));
    OR4 OR4_156 (.A(OR4_570_Y), .B(OR2_77_Y), .C(
        \Z\R_DATA_TEMPR22[42] ), .D(\Z\R_DATA_TEMPR23[42] ), .Y(
        OR4_156_Y));
    OR4 OR4_535 (.A(\Z\R_DATA_TEMPR24[15] ), .B(\Z\R_DATA_TEMPR25[15] )
        , .C(\Z\R_DATA_TEMPR26[15] ), .D(\Z\R_DATA_TEMPR27[15] ), .Y(
        OR4_535_Y));
    OR2 OR2_36 (.A(\Z\R_DATA_TEMPR20[34] ), .B(\Z\R_DATA_TEMPR21[34] ), 
        .Y(OR2_36_Y));
    OR4 OR4_68 (.A(\Z\R_DATA_TEMPR24[26] ), .B(\Z\R_DATA_TEMPR25[26] ), 
        .C(\Z\R_DATA_TEMPR26[26] ), .D(\Z\R_DATA_TEMPR27[26] ), .Y(
        OR4_68_Y));
    OR2 OR2_24 (.A(\Z\R_DATA_TEMPR20[23] ), .B(\Z\R_DATA_TEMPR21[23] ), 
        .Y(OR2_24_Y));
    OR4 OR4_377 (.A(\Z\R_DATA_TEMPR16[38] ), .B(\Z\R_DATA_TEMPR17[38] )
        , .C(\Z\R_DATA_TEMPR18[38] ), .D(\Z\R_DATA_TEMPR19[38] ), .Y(
        OR4_377_Y));
    OR4 OR4_170 (.A(OR4_415_Y), .B(OR4_540_Y), .C(OR4_538_Y), .D(
        OR4_653_Y), .Y(OR4_170_Y));
    OR4 OR4_708 (.A(OR4_175_Y), .B(OR2_26_Y), .C(
        \Z\R_DATA_TEMPR22[54] ), .D(\Z\R_DATA_TEMPR23[54] ), .Y(
        OR4_708_Y));
    OR4 OR4_626 (.A(\Z\R_DATA_TEMPR0[72] ), .B(\Z\R_DATA_TEMPR1[72] ), 
        .C(\Z\R_DATA_TEMPR2[72] ), .D(\Z\R_DATA_TEMPR3[72] ), .Y(
        OR4_626_Y));
    OR4 OR4_31 (.A(\Z\R_DATA_TEMPR4[63] ), .B(\Z\R_DATA_TEMPR5[63] ), 
        .C(\Z\R_DATA_TEMPR6[63] ), .D(\Z\R_DATA_TEMPR7[63] ), .Y(
        OR4_31_Y));
    OR4 \OR4_R_DATA[65]  (.A(OR4_115_Y), .B(OR4_468_Y), .C(OR4_28_Y), 
        .D(OR4_546_Y), .Y(R_DATA_c[65]));
    OR4 OR4_633 (.A(OR4_405_Y), .B(OR4_268_Y), .C(OR4_132_Y), .D(
        OR4_172_Y), .Y(OR4_633_Y));
    OR4 \OR4_R_DATA[31]  (.A(OR4_170_Y), .B(OR4_126_Y), .C(OR4_142_Y), 
        .D(OR4_648_Y), .Y(R_DATA_c[31]));
    OR4 OR4_385 (.A(\Z\R_DATA_TEMPR8[67] ), .B(\Z\R_DATA_TEMPR9[67] ), 
        .C(\Z\R_DATA_TEMPR10[67] ), .D(\Z\R_DATA_TEMPR11[67] ), .Y(
        OR4_385_Y));
    OR4 OR4_243 (.A(\Z\R_DATA_TEMPR24[34] ), .B(\Z\R_DATA_TEMPR25[34] )
        , .C(\Z\R_DATA_TEMPR26[34] ), .D(\Z\R_DATA_TEMPR27[34] ), .Y(
        OR4_243_Y));
    OR4 OR4_394 (.A(\Z\R_DATA_TEMPR16[61] ), .B(\Z\R_DATA_TEMPR17[61] )
        , .C(\Z\R_DATA_TEMPR18[61] ), .D(\Z\R_DATA_TEMPR19[61] ), .Y(
        OR4_394_Y));
    OR4 OR4_358 (.A(OR4_490_Y), .B(OR2_46_Y), .C(\Z\R_DATA_TEMPR22[2] )
        , .D(\Z\R_DATA_TEMPR23[2] ), .Y(OR4_358_Y));
    OR4 OR4_80 (.A(\Z\R_DATA_TEMPR12[22] ), .B(\Z\R_DATA_TEMPR13[22] ), 
        .C(\Z\R_DATA_TEMPR14[22] ), .D(\Z\R_DATA_TEMPR15[22] ), .Y(
        OR4_80_Y));
    OR4 OR4_191 (.A(OR4_683_Y), .B(OR4_537_Y), .C(OR4_413_Y), .D(
        OR4_444_Y), .Y(OR4_191_Y));
    OR4 OR4_108 (.A(\Z\R_DATA_TEMPR12[72] ), .B(\Z\R_DATA_TEMPR13[72] )
        , .C(\Z\R_DATA_TEMPR14[72] ), .D(\Z\R_DATA_TEMPR15[72] ), .Y(
        OR4_108_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%12%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C1 (
        .A_DOUT({\Z\R_DATA_TEMPR12[79] , \Z\R_DATA_TEMPR12[78] , 
        \Z\R_DATA_TEMPR12[77] , \Z\R_DATA_TEMPR12[76] , 
        \Z\R_DATA_TEMPR12[75] , \Z\R_DATA_TEMPR12[74] , 
        \Z\R_DATA_TEMPR12[73] , \Z\R_DATA_TEMPR12[72] , 
        \Z\R_DATA_TEMPR12[71] , \Z\R_DATA_TEMPR12[70] , 
        \Z\R_DATA_TEMPR12[69] , \Z\R_DATA_TEMPR12[68] , 
        \Z\R_DATA_TEMPR12[67] , \Z\R_DATA_TEMPR12[66] , 
        \Z\R_DATA_TEMPR12[65] , \Z\R_DATA_TEMPR12[64] , 
        \Z\R_DATA_TEMPR12[63] , \Z\R_DATA_TEMPR12[62] , 
        \Z\R_DATA_TEMPR12[61] , \Z\R_DATA_TEMPR12[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR12[59] , \Z\R_DATA_TEMPR12[58] , 
        \Z\R_DATA_TEMPR12[57] , \Z\R_DATA_TEMPR12[56] , 
        \Z\R_DATA_TEMPR12[55] , \Z\R_DATA_TEMPR12[54] , 
        \Z\R_DATA_TEMPR12[53] , \Z\R_DATA_TEMPR12[52] , 
        \Z\R_DATA_TEMPR12[51] , \Z\R_DATA_TEMPR12[50] , 
        \Z\R_DATA_TEMPR12[49] , \Z\R_DATA_TEMPR12[48] , 
        \Z\R_DATA_TEMPR12[47] , \Z\R_DATA_TEMPR12[46] , 
        \Z\R_DATA_TEMPR12[45] , \Z\R_DATA_TEMPR12[44] , 
        \Z\R_DATA_TEMPR12[43] , \Z\R_DATA_TEMPR12[42] , 
        \Z\R_DATA_TEMPR12[41] , \Z\R_DATA_TEMPR12[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[12][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[3] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[3] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_1 (.A(\Z\R_DATA_TEMPR8[66] ), .B(\Z\R_DATA_TEMPR9[66] ), 
        .C(\Z\R_DATA_TEMPR10[66] ), .D(\Z\R_DATA_TEMPR11[66] ), .Y(
        OR4_1_Y));
    OR2 OR2_40 (.A(\Z\R_DATA_TEMPR20[20] ), .B(\Z\R_DATA_TEMPR21[20] ), 
        .Y(OR2_40_Y));
    OR4 OR4_87 (.A(OR4_151_Y), .B(OR4_554_Y), .C(OR4_98_Y), .D(
        OR4_450_Y), .Y(OR4_87_Y));
    OR4 \OR4_R_DATA[30]  (.A(OR4_37_Y), .B(OR4_214_Y), .C(OR4_529_Y), 
        .D(OR4_264_Y), .Y(R_DATA_c[30]));
    OR4 OR4_178 (.A(OR4_224_Y), .B(OR4_453_Y), .C(OR4_642_Y), .D(
        OR4_254_Y), .Y(OR4_178_Y));
    OR2 OR2_47 (.A(\Z\R_DATA_TEMPR20[17] ), .B(\Z\R_DATA_TEMPR21[17] ), 
        .Y(OR2_47_Y));
    OR4 OR4_159 (.A(\Z\R_DATA_TEMPR8[42] ), .B(\Z\R_DATA_TEMPR9[42] ), 
        .C(\Z\R_DATA_TEMPR10[42] ), .D(\Z\R_DATA_TEMPR11[42] ), .Y(
        OR4_159_Y));
    OR4 OR4_491 (.A(\Z\R_DATA_TEMPR12[11] ), .B(\Z\R_DATA_TEMPR13[11] )
        , .C(\Z\R_DATA_TEMPR14[11] ), .D(\Z\R_DATA_TEMPR15[11] ), .Y(
        OR4_491_Y));
    OR4 OR4_165 (.A(\Z\R_DATA_TEMPR16[72] ), .B(\Z\R_DATA_TEMPR17[72] )
        , .C(\Z\R_DATA_TEMPR18[72] ), .D(\Z\R_DATA_TEMPR19[72] ), .Y(
        OR4_165_Y));
    OR4 OR4_133 (.A(OR4_483_Y), .B(OR2_27_Y), .C(
        \Z\R_DATA_TEMPR22[58] ), .D(\Z\R_DATA_TEMPR23[58] ), .Y(
        OR4_133_Y));
    OR4 OR4_515 (.A(OR4_140_Y), .B(OR2_19_Y), .C(\Z\R_DATA_TEMPR22[6] )
        , .D(\Z\R_DATA_TEMPR23[6] ), .Y(OR4_515_Y));
    OR4 OR4_498 (.A(\Z\R_DATA_TEMPR8[73] ), .B(\Z\R_DATA_TEMPR9[73] ), 
        .C(\Z\R_DATA_TEMPR10[73] ), .D(\Z\R_DATA_TEMPR11[73] ), .Y(
        OR4_498_Y));
    OR4 \OR4_R_DATA[36]  (.A(OR4_504_Y), .B(OR4_176_Y), .C(OR4_302_Y), 
        .D(OR4_332_Y), .Y(R_DATA_c[36]));
    OR4 OR4_92 (.A(\Z\R_DATA_TEMPR0[6] ), .B(\Z\R_DATA_TEMPR1[6] ), .C(
        \Z\R_DATA_TEMPR2[6] ), .D(\Z\R_DATA_TEMPR3[6] ), .Y(OR4_92_Y));
    OR4 OR4_467 (.A(\Z\R_DATA_TEMPR0[18] ), .B(\Z\R_DATA_TEMPR1[18] ), 
        .C(\Z\R_DATA_TEMPR2[18] ), .D(\Z\R_DATA_TEMPR3[18] ), .Y(
        OR4_467_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[1]  (.A(CFG2_6_Y), .B(
        R_ADDR_c[13]), .C(R_EN_c), .Y(\Z\BLKY2[1] ));
    OR4 OR4_648 (.A(\Z\R_DATA_TEMPR28[31] ), .B(\Z\R_DATA_TEMPR29[31] )
        , .C(\Z\R_DATA_TEMPR30[31] ), .D(\Z\R_DATA_TEMPR31[31] ), .Y(
        OR4_648_Y));
    OR4 OR4_685 (.A(\Z\R_DATA_TEMPR0[39] ), .B(\Z\R_DATA_TEMPR1[39] ), 
        .C(\Z\R_DATA_TEMPR2[39] ), .D(\Z\R_DATA_TEMPR3[39] ), .Y(
        OR4_685_Y));
    OR2 OR2_60 (.A(\Z\R_DATA_TEMPR20[64] ), .B(\Z\R_DATA_TEMPR21[64] ), 
        .Y(OR2_60_Y));
    OR4 OR4_613 (.A(\Z\R_DATA_TEMPR12[76] ), .B(\Z\R_DATA_TEMPR13[76] )
        , .C(\Z\R_DATA_TEMPR14[76] ), .D(\Z\R_DATA_TEMPR15[76] ), .Y(
        OR4_613_Y));
    OR2 OR2_74 (.A(\Z\R_DATA_TEMPR20[36] ), .B(\Z\R_DATA_TEMPR21[36] ), 
        .Y(OR2_74_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%26%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0 (
        .A_DOUT({\Z\R_DATA_TEMPR26[39] , \Z\R_DATA_TEMPR26[38] , 
        \Z\R_DATA_TEMPR26[37] , \Z\R_DATA_TEMPR26[36] , 
        \Z\R_DATA_TEMPR26[35] , \Z\R_DATA_TEMPR26[34] , 
        \Z\R_DATA_TEMPR26[33] , \Z\R_DATA_TEMPR26[32] , 
        \Z\R_DATA_TEMPR26[31] , \Z\R_DATA_TEMPR26[30] , 
        \Z\R_DATA_TEMPR26[29] , \Z\R_DATA_TEMPR26[28] , 
        \Z\R_DATA_TEMPR26[27] , \Z\R_DATA_TEMPR26[26] , 
        \Z\R_DATA_TEMPR26[25] , \Z\R_DATA_TEMPR26[24] , 
        \Z\R_DATA_TEMPR26[23] , \Z\R_DATA_TEMPR26[22] , 
        \Z\R_DATA_TEMPR26[21] , \Z\R_DATA_TEMPR26[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR26[19] , \Z\R_DATA_TEMPR26[18] , 
        \Z\R_DATA_TEMPR26[17] , \Z\R_DATA_TEMPR26[16] , 
        \Z\R_DATA_TEMPR26[15] , \Z\R_DATA_TEMPR26[14] , 
        \Z\R_DATA_TEMPR26[13] , \Z\R_DATA_TEMPR26[12] , 
        \Z\R_DATA_TEMPR26[11] , \Z\R_DATA_TEMPR26[10] , 
        \Z\R_DATA_TEMPR26[9] , \Z\R_DATA_TEMPR26[8] , 
        \Z\R_DATA_TEMPR26[7] , \Z\R_DATA_TEMPR26[6] , 
        \Z\R_DATA_TEMPR26[5] , \Z\R_DATA_TEMPR26[4] , 
        \Z\R_DATA_TEMPR26[3] , \Z\R_DATA_TEMPR26[2] , 
        \Z\R_DATA_TEMPR26[1] , \Z\R_DATA_TEMPR26[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[26][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[6] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[6] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_642 (.A(\Z\R_DATA_TEMPR8[3] ), .B(\Z\R_DATA_TEMPR9[3] ), 
        .C(\Z\R_DATA_TEMPR10[3] ), .D(\Z\R_DATA_TEMPR11[3] ), .Y(
        OR4_642_Y));
    OR2 OR2_67 (.A(\Z\R_DATA_TEMPR20[16] ), .B(\Z\R_DATA_TEMPR21[16] ), 
        .Y(OR2_67_Y));
    OR2 OR2_30 (.A(\Z\R_DATA_TEMPR20[35] ), .B(\Z\R_DATA_TEMPR21[35] ), 
        .Y(OR2_30_Y));
    CFG2 #( .INIT(4'h8) )  CFG2_0 (.A(W_ADDR_c[12]), .B(W_ADDR_c[11]), 
        .Y(CFG2_0_Y));
    OR4 OR4_324 (.A(\Z\R_DATA_TEMPR24[54] ), .B(\Z\R_DATA_TEMPR25[54] )
        , .C(\Z\R_DATA_TEMPR26[54] ), .D(\Z\R_DATA_TEMPR27[54] ), .Y(
        OR4_324_Y));
    OR4 OR4_265 (.A(OR4_695_Y), .B(OR2_18_Y), .C(
        \Z\R_DATA_TEMPR22[15] ), .D(\Z\R_DATA_TEMPR23[15] ), .Y(
        OR4_265_Y));
    OR4 OR4_49 (.A(\Z\R_DATA_TEMPR24[42] ), .B(\Z\R_DATA_TEMPR25[42] ), 
        .C(\Z\R_DATA_TEMPR26[42] ), .D(\Z\R_DATA_TEMPR27[42] ), .Y(
        OR4_49_Y));
    OR4 OR4_599 (.A(OR4_573_Y), .B(OR4_568_Y), .C(OR4_525_Y), .D(
        OR4_702_Y), .Y(OR4_599_Y));
    OR2 OR2_14 (.A(\Z\R_DATA_TEMPR20[32] ), .B(\Z\R_DATA_TEMPR21[32] ), 
        .Y(OR2_14_Y));
    OR2 OR2_37 (.A(\Z\R_DATA_TEMPR20[38] ), .B(\Z\R_DATA_TEMPR21[38] ), 
        .Y(OR2_37_Y));
    OR4 OR4_590 (.A(\Z\R_DATA_TEMPR4[61] ), .B(\Z\R_DATA_TEMPR5[61] ), 
        .C(\Z\R_DATA_TEMPR6[61] ), .D(\Z\R_DATA_TEMPR7[61] ), .Y(
        OR4_590_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%30%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0 (
        .A_DOUT({\Z\R_DATA_TEMPR30[39] , \Z\R_DATA_TEMPR30[38] , 
        \Z\R_DATA_TEMPR30[37] , \Z\R_DATA_TEMPR30[36] , 
        \Z\R_DATA_TEMPR30[35] , \Z\R_DATA_TEMPR30[34] , 
        \Z\R_DATA_TEMPR30[33] , \Z\R_DATA_TEMPR30[32] , 
        \Z\R_DATA_TEMPR30[31] , \Z\R_DATA_TEMPR30[30] , 
        \Z\R_DATA_TEMPR30[29] , \Z\R_DATA_TEMPR30[28] , 
        \Z\R_DATA_TEMPR30[27] , \Z\R_DATA_TEMPR30[26] , 
        \Z\R_DATA_TEMPR30[25] , \Z\R_DATA_TEMPR30[24] , 
        \Z\R_DATA_TEMPR30[23] , \Z\R_DATA_TEMPR30[22] , 
        \Z\R_DATA_TEMPR30[21] , \Z\R_DATA_TEMPR30[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR30[19] , \Z\R_DATA_TEMPR30[18] , 
        \Z\R_DATA_TEMPR30[17] , \Z\R_DATA_TEMPR30[16] , 
        \Z\R_DATA_TEMPR30[15] , \Z\R_DATA_TEMPR30[14] , 
        \Z\R_DATA_TEMPR30[13] , \Z\R_DATA_TEMPR30[12] , 
        \Z\R_DATA_TEMPR30[11] , \Z\R_DATA_TEMPR30[10] , 
        \Z\R_DATA_TEMPR30[9] , \Z\R_DATA_TEMPR30[8] , 
        \Z\R_DATA_TEMPR30[7] , \Z\R_DATA_TEMPR30[6] , 
        \Z\R_DATA_TEMPR30[5] , \Z\R_DATA_TEMPR30[4] , 
        \Z\R_DATA_TEMPR30[3] , \Z\R_DATA_TEMPR30[2] , 
        \Z\R_DATA_TEMPR30[1] , \Z\R_DATA_TEMPR30[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[30][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[7] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[7] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_121 (.A(\Z\R_DATA_TEMPR0[36] ), .B(\Z\R_DATA_TEMPR1[36] ), 
        .C(\Z\R_DATA_TEMPR2[36] ), .D(\Z\R_DATA_TEMPR3[36] ), .Y(
        OR4_121_Y));
    OR2 OR2_53 (.A(\Z\R_DATA_TEMPR20[65] ), .B(\Z\R_DATA_TEMPR21[65] ), 
        .Y(OR2_53_Y));
    OR4 \OR4_R_DATA[18]  (.A(OR4_689_Y), .B(OR4_594_Y), .C(OR4_272_Y), 
        .D(OR4_361_Y), .Y(R_DATA_c[18]));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%3%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C1 (
        .A_DOUT({\Z\R_DATA_TEMPR3[79] , \Z\R_DATA_TEMPR3[78] , 
        \Z\R_DATA_TEMPR3[77] , \Z\R_DATA_TEMPR3[76] , 
        \Z\R_DATA_TEMPR3[75] , \Z\R_DATA_TEMPR3[74] , 
        \Z\R_DATA_TEMPR3[73] , \Z\R_DATA_TEMPR3[72] , 
        \Z\R_DATA_TEMPR3[71] , \Z\R_DATA_TEMPR3[70] , 
        \Z\R_DATA_TEMPR3[69] , \Z\R_DATA_TEMPR3[68] , 
        \Z\R_DATA_TEMPR3[67] , \Z\R_DATA_TEMPR3[66] , 
        \Z\R_DATA_TEMPR3[65] , \Z\R_DATA_TEMPR3[64] , 
        \Z\R_DATA_TEMPR3[63] , \Z\R_DATA_TEMPR3[62] , 
        \Z\R_DATA_TEMPR3[61] , \Z\R_DATA_TEMPR3[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR3[59] , \Z\R_DATA_TEMPR3[58] , 
        \Z\R_DATA_TEMPR3[57] , \Z\R_DATA_TEMPR3[56] , 
        \Z\R_DATA_TEMPR3[55] , \Z\R_DATA_TEMPR3[54] , 
        \Z\R_DATA_TEMPR3[53] , \Z\R_DATA_TEMPR3[52] , 
        \Z\R_DATA_TEMPR3[51] , \Z\R_DATA_TEMPR3[50] , 
        \Z\R_DATA_TEMPR3[49] , \Z\R_DATA_TEMPR3[48] , 
        \Z\R_DATA_TEMPR3[47] , \Z\R_DATA_TEMPR3[46] , 
        \Z\R_DATA_TEMPR3[45] , \Z\R_DATA_TEMPR3[44] , 
        \Z\R_DATA_TEMPR3[43] , \Z\R_DATA_TEMPR3[42] , 
        \Z\R_DATA_TEMPR3[41] , \Z\R_DATA_TEMPR3[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[3][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[0] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[0] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%1%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C1 (
        .A_DOUT({\Z\R_DATA_TEMPR1[79] , \Z\R_DATA_TEMPR1[78] , 
        \Z\R_DATA_TEMPR1[77] , \Z\R_DATA_TEMPR1[76] , 
        \Z\R_DATA_TEMPR1[75] , \Z\R_DATA_TEMPR1[74] , 
        \Z\R_DATA_TEMPR1[73] , \Z\R_DATA_TEMPR1[72] , 
        \Z\R_DATA_TEMPR1[71] , \Z\R_DATA_TEMPR1[70] , 
        \Z\R_DATA_TEMPR1[69] , \Z\R_DATA_TEMPR1[68] , 
        \Z\R_DATA_TEMPR1[67] , \Z\R_DATA_TEMPR1[66] , 
        \Z\R_DATA_TEMPR1[65] , \Z\R_DATA_TEMPR1[64] , 
        \Z\R_DATA_TEMPR1[63] , \Z\R_DATA_TEMPR1[62] , 
        \Z\R_DATA_TEMPR1[61] , \Z\R_DATA_TEMPR1[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR1[59] , \Z\R_DATA_TEMPR1[58] , 
        \Z\R_DATA_TEMPR1[57] , \Z\R_DATA_TEMPR1[56] , 
        \Z\R_DATA_TEMPR1[55] , \Z\R_DATA_TEMPR1[54] , 
        \Z\R_DATA_TEMPR1[53] , \Z\R_DATA_TEMPR1[52] , 
        \Z\R_DATA_TEMPR1[51] , \Z\R_DATA_TEMPR1[50] , 
        \Z\R_DATA_TEMPR1[49] , \Z\R_DATA_TEMPR1[48] , 
        \Z\R_DATA_TEMPR1[47] , \Z\R_DATA_TEMPR1[46] , 
        \Z\R_DATA_TEMPR1[45] , \Z\R_DATA_TEMPR1[44] , 
        \Z\R_DATA_TEMPR1[43] , \Z\R_DATA_TEMPR1[42] , 
        \Z\R_DATA_TEMPR1[41] , \Z\R_DATA_TEMPR1[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[1][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[0] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[0] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_680 (.A(OR4_99_Y), .B(OR2_69_Y), .C(\Z\R_DATA_TEMPR22[0] ), 
        .D(\Z\R_DATA_TEMPR23[0] ), .Y(OR4_680_Y));
    OR4 OR4_132 (.A(\Z\R_DATA_TEMPR8[28] ), .B(\Z\R_DATA_TEMPR9[28] ), 
        .C(\Z\R_DATA_TEMPR10[28] ), .D(\Z\R_DATA_TEMPR11[28] ), .Y(
        OR4_132_Y));
    OR4 OR4_113 (.A(\Z\R_DATA_TEMPR16[13] ), .B(\Z\R_DATA_TEMPR17[13] )
        , .C(\Z\R_DATA_TEMPR18[13] ), .D(\Z\R_DATA_TEMPR19[13] ), .Y(
        OR4_113_Y));
    OR4 OR4_7 (.A(\Z\R_DATA_TEMPR4[79] ), .B(\Z\R_DATA_TEMPR5[79] ), 
        .C(\Z\R_DATA_TEMPR6[79] ), .D(\Z\R_DATA_TEMPR7[79] ), .Y(
        OR4_7_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%11%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C1 (
        .A_DOUT({\Z\R_DATA_TEMPR11[79] , \Z\R_DATA_TEMPR11[78] , 
        \Z\R_DATA_TEMPR11[77] , \Z\R_DATA_TEMPR11[76] , 
        \Z\R_DATA_TEMPR11[75] , \Z\R_DATA_TEMPR11[74] , 
        \Z\R_DATA_TEMPR11[73] , \Z\R_DATA_TEMPR11[72] , 
        \Z\R_DATA_TEMPR11[71] , \Z\R_DATA_TEMPR11[70] , 
        \Z\R_DATA_TEMPR11[69] , \Z\R_DATA_TEMPR11[68] , 
        \Z\R_DATA_TEMPR11[67] , \Z\R_DATA_TEMPR11[66] , 
        \Z\R_DATA_TEMPR11[65] , \Z\R_DATA_TEMPR11[64] , 
        \Z\R_DATA_TEMPR11[63] , \Z\R_DATA_TEMPR11[62] , 
        \Z\R_DATA_TEMPR11[61] , \Z\R_DATA_TEMPR11[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR11[59] , \Z\R_DATA_TEMPR11[58] , 
        \Z\R_DATA_TEMPR11[57] , \Z\R_DATA_TEMPR11[56] , 
        \Z\R_DATA_TEMPR11[55] , \Z\R_DATA_TEMPR11[54] , 
        \Z\R_DATA_TEMPR11[53] , \Z\R_DATA_TEMPR11[52] , 
        \Z\R_DATA_TEMPR11[51] , \Z\R_DATA_TEMPR11[50] , 
        \Z\R_DATA_TEMPR11[49] , \Z\R_DATA_TEMPR11[48] , 
        \Z\R_DATA_TEMPR11[47] , \Z\R_DATA_TEMPR11[46] , 
        \Z\R_DATA_TEMPR11[45] , \Z\R_DATA_TEMPR11[44] , 
        \Z\R_DATA_TEMPR11[43] , \Z\R_DATA_TEMPR11[42] , 
        \Z\R_DATA_TEMPR11[41] , \Z\R_DATA_TEMPR11[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[11][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[2] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[2] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_421 (.A(OR4_484_Y), .B(OR4_158_Y), .C(OR4_429_Y), .D(
        OR4_55_Y), .Y(OR4_421_Y));
    OR4 OR4_463 (.A(\Z\R_DATA_TEMPR12[4] ), .B(\Z\R_DATA_TEMPR13[4] ), 
        .C(\Z\R_DATA_TEMPR14[4] ), .D(\Z\R_DATA_TEMPR15[4] ), .Y(
        OR4_463_Y));
    OR4 OR4_661 (.A(OR4_211_Y), .B(OR2_49_Y), .C(\Z\R_DATA_TEMPR22[7] )
        , .D(\Z\R_DATA_TEMPR23[7] ), .Y(OR4_661_Y));
    OR4 OR4_657 (.A(\Z\R_DATA_TEMPR24[77] ), .B(\Z\R_DATA_TEMPR25[77] )
        , .C(\Z\R_DATA_TEMPR26[77] ), .D(\Z\R_DATA_TEMPR27[77] ), .Y(
        OR4_657_Y));
    OR4 OR4_428 (.A(OR4_631_Y), .B(OR2_28_Y), .C(
        \Z\R_DATA_TEMPR22[14] ), .D(\Z\R_DATA_TEMPR23[14] ), .Y(
        OR4_428_Y));
    OR4 OR4_268 (.A(\Z\R_DATA_TEMPR4[28] ), .B(\Z\R_DATA_TEMPR5[28] ), 
        .C(\Z\R_DATA_TEMPR6[28] ), .D(\Z\R_DATA_TEMPR7[28] ), .Y(
        OR4_268_Y));
    OR4 OR4_387 (.A(\Z\R_DATA_TEMPR8[8] ), .B(\Z\R_DATA_TEMPR9[8] ), 
        .C(\Z\R_DATA_TEMPR10[8] ), .D(\Z\R_DATA_TEMPR11[8] ), .Y(
        OR4_387_Y));
    OR4 OR4_180 (.A(\Z\R_DATA_TEMPR28[73] ), .B(\Z\R_DATA_TEMPR29[73] )
        , .C(\Z\R_DATA_TEMPR30[73] ), .D(\Z\R_DATA_TEMPR31[73] ), .Y(
        OR4_180_Y));
    OR4 OR4_105 (.A(\Z\R_DATA_TEMPR16[5] ), .B(\Z\R_DATA_TEMPR17[5] ), 
        .C(\Z\R_DATA_TEMPR18[5] ), .D(\Z\R_DATA_TEMPR19[5] ), .Y(
        OR4_105_Y));
    OR4 OR4_407 (.A(\Z\R_DATA_TEMPR4[26] ), .B(\Z\R_DATA_TEMPR5[26] ), 
        .C(\Z\R_DATA_TEMPR6[26] ), .D(\Z\R_DATA_TEMPR7[26] ), .Y(
        OR4_407_Y));
    OR4 OR4_393 (.A(OR4_685_Y), .B(OR4_221_Y), .C(OR4_519_Y), .D(
        OR4_85_Y), .Y(OR4_393_Y));
    OR4 OR4_175 (.A(\Z\R_DATA_TEMPR16[54] ), .B(\Z\R_DATA_TEMPR17[54] )
        , .C(\Z\R_DATA_TEMPR18[54] ), .D(\Z\R_DATA_TEMPR19[54] ), .Y(
        OR4_175_Y));
    OR4 OR4_239 (.A(\Z\R_DATA_TEMPR0[9] ), .B(\Z\R_DATA_TEMPR1[9] ), 
        .C(\Z\R_DATA_TEMPR2[9] ), .D(\Z\R_DATA_TEMPR3[9] ), .Y(
        OR4_239_Y));
    OR4 OR4_42 (.A(OR4_357_Y), .B(OR2_33_Y), .C(\Z\R_DATA_TEMPR22[79] )
        , .D(\Z\R_DATA_TEMPR23[79] ), .Y(OR4_42_Y));
    OR4 OR4_529 (.A(\Z\R_DATA_TEMPR24[30] ), .B(\Z\R_DATA_TEMPR25[30] )
        , .C(\Z\R_DATA_TEMPR26[30] ), .D(\Z\R_DATA_TEMPR27[30] ), .Y(
        OR4_529_Y));
    OR4 OR4_477 (.A(\Z\R_DATA_TEMPR4[23] ), .B(\Z\R_DATA_TEMPR5[23] ), 
        .C(\Z\R_DATA_TEMPR6[23] ), .D(\Z\R_DATA_TEMPR7[23] ), .Y(
        OR4_477_Y));
    OR4 OR4_492 (.A(\Z\R_DATA_TEMPR0[79] ), .B(\Z\R_DATA_TEMPR1[79] ), 
        .C(\Z\R_DATA_TEMPR2[79] ), .D(\Z\R_DATA_TEMPR3[79] ), .Y(
        OR4_492_Y));
    OR4 OR4_520 (.A(OR4_251_Y), .B(OR2_17_Y), .C(
        \Z\R_DATA_TEMPR22[55] ), .D(\Z\R_DATA_TEMPR23[55] ), .Y(
        OR4_520_Y));
    OR2 OR2_51 (.A(\Z\R_DATA_TEMPR20[24] ), .B(\Z\R_DATA_TEMPR21[24] ), 
        .Y(OR2_51_Y));
    OR4 OR4_88 (.A(OR4_325_Y), .B(OR4_201_Y), .C(OR4_185_Y), .D(
        OR4_620_Y), .Y(OR4_88_Y));
    OR4 OR4_499 (.A(\Z\R_DATA_TEMPR24[2] ), .B(\Z\R_DATA_TEMPR25[2] ), 
        .C(\Z\R_DATA_TEMPR26[2] ), .D(\Z\R_DATA_TEMPR27[2] ), .Y(
        OR4_499_Y));
    OR4 OR4_205 (.A(OR4_637_Y), .B(OR2_44_Y), .C(
        \Z\R_DATA_TEMPR22[25] ), .D(\Z\R_DATA_TEMPR23[25] ), .Y(
        OR4_205_Y));
    OR4 OR4_188 (.A(\Z\R_DATA_TEMPR0[66] ), .B(\Z\R_DATA_TEMPR1[66] ), 
        .C(\Z\R_DATA_TEMPR2[66] ), .D(\Z\R_DATA_TEMPR3[66] ), .Y(
        OR4_188_Y));
    OR4 OR4_196 (.A(\Z\R_DATA_TEMPR8[55] ), .B(\Z\R_DATA_TEMPR9[55] ), 
        .C(\Z\R_DATA_TEMPR10[55] ), .D(\Z\R_DATA_TEMPR11[55] ), .Y(
        OR4_196_Y));
    OR4 OR4_112 (.A(\Z\R_DATA_TEMPR16[64] ), .B(\Z\R_DATA_TEMPR17[64] )
        , .C(\Z\R_DATA_TEMPR18[64] ), .D(\Z\R_DATA_TEMPR19[64] ), .Y(
        OR4_112_Y));
    OR2 OR2_48 (.A(\Z\R_DATA_TEMPR20[49] ), .B(\Z\R_DATA_TEMPR21[49] ), 
        .Y(OR2_48_Y));
    OR4 \OR4_R_DATA[48]  (.A(OR4_338_Y), .B(OR4_258_Y), .C(OR4_641_Y), 
        .D(OR4_13_Y), .Y(R_DATA_c[48]));
    OR4 OR4_275 (.A(\Z\R_DATA_TEMPR24[8] ), .B(\Z\R_DATA_TEMPR25[8] ), 
        .C(\Z\R_DATA_TEMPR26[8] ), .D(\Z\R_DATA_TEMPR27[8] ), .Y(
        OR4_275_Y));
    OR4 OR4_646 (.A(\Z\R_DATA_TEMPR8[15] ), .B(\Z\R_DATA_TEMPR9[15] ), 
        .C(\Z\R_DATA_TEMPR10[15] ), .D(\Z\R_DATA_TEMPR11[15] ), .Y(
        OR4_646_Y));
    OR4 \OR4_R_DATA[37]  (.A(OR4_316_Y), .B(OR4_670_Y), .C(OR4_119_Y), 
        .D(OR4_208_Y), .Y(R_DATA_c[37]));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%25%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C1 (
        .A_DOUT({\Z\R_DATA_TEMPR25[79] , \Z\R_DATA_TEMPR25[78] , 
        \Z\R_DATA_TEMPR25[77] , \Z\R_DATA_TEMPR25[76] , 
        \Z\R_DATA_TEMPR25[75] , \Z\R_DATA_TEMPR25[74] , 
        \Z\R_DATA_TEMPR25[73] , \Z\R_DATA_TEMPR25[72] , 
        \Z\R_DATA_TEMPR25[71] , \Z\R_DATA_TEMPR25[70] , 
        \Z\R_DATA_TEMPR25[69] , \Z\R_DATA_TEMPR25[68] , 
        \Z\R_DATA_TEMPR25[67] , \Z\R_DATA_TEMPR25[66] , 
        \Z\R_DATA_TEMPR25[65] , \Z\R_DATA_TEMPR25[64] , 
        \Z\R_DATA_TEMPR25[63] , \Z\R_DATA_TEMPR25[62] , 
        \Z\R_DATA_TEMPR25[61] , \Z\R_DATA_TEMPR25[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR25[59] , \Z\R_DATA_TEMPR25[58] , 
        \Z\R_DATA_TEMPR25[57] , \Z\R_DATA_TEMPR25[56] , 
        \Z\R_DATA_TEMPR25[55] , \Z\R_DATA_TEMPR25[54] , 
        \Z\R_DATA_TEMPR25[53] , \Z\R_DATA_TEMPR25[52] , 
        \Z\R_DATA_TEMPR25[51] , \Z\R_DATA_TEMPR25[50] , 
        \Z\R_DATA_TEMPR25[49] , \Z\R_DATA_TEMPR25[48] , 
        \Z\R_DATA_TEMPR25[47] , \Z\R_DATA_TEMPR25[46] , 
        \Z\R_DATA_TEMPR25[45] , \Z\R_DATA_TEMPR25[44] , 
        \Z\R_DATA_TEMPR25[43] , \Z\R_DATA_TEMPR25[42] , 
        \Z\R_DATA_TEMPR25[41] , \Z\R_DATA_TEMPR25[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[25][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[6] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[6] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_257 (.A(\Z\R_DATA_TEMPR28[67] ), .B(\Z\R_DATA_TEMPR29[67] )
        , .C(\Z\R_DATA_TEMPR30[67] ), .D(\Z\R_DATA_TEMPR31[67] ), .Y(
        OR4_257_Y));
    OR4 OR4_398 (.A(\Z\R_DATA_TEMPR24[12] ), .B(\Z\R_DATA_TEMPR25[12] )
        , .C(\Z\R_DATA_TEMPR26[12] ), .D(\Z\R_DATA_TEMPR27[12] ), .Y(
        OR4_398_Y));
    OR4 OR4_157 (.A(\Z\R_DATA_TEMPR12[9] ), .B(\Z\R_DATA_TEMPR13[9] ), 
        .C(\Z\R_DATA_TEMPR14[9] ), .D(\Z\R_DATA_TEMPR15[9] ), .Y(
        OR4_157_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%5%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C1 (
        .A_DOUT({\Z\R_DATA_TEMPR5[79] , \Z\R_DATA_TEMPR5[78] , 
        \Z\R_DATA_TEMPR5[77] , \Z\R_DATA_TEMPR5[76] , 
        \Z\R_DATA_TEMPR5[75] , \Z\R_DATA_TEMPR5[74] , 
        \Z\R_DATA_TEMPR5[73] , \Z\R_DATA_TEMPR5[72] , 
        \Z\R_DATA_TEMPR5[71] , \Z\R_DATA_TEMPR5[70] , 
        \Z\R_DATA_TEMPR5[69] , \Z\R_DATA_TEMPR5[68] , 
        \Z\R_DATA_TEMPR5[67] , \Z\R_DATA_TEMPR5[66] , 
        \Z\R_DATA_TEMPR5[65] , \Z\R_DATA_TEMPR5[64] , 
        \Z\R_DATA_TEMPR5[63] , \Z\R_DATA_TEMPR5[62] , 
        \Z\R_DATA_TEMPR5[61] , \Z\R_DATA_TEMPR5[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR5[59] , \Z\R_DATA_TEMPR5[58] , 
        \Z\R_DATA_TEMPR5[57] , \Z\R_DATA_TEMPR5[56] , 
        \Z\R_DATA_TEMPR5[55] , \Z\R_DATA_TEMPR5[54] , 
        \Z\R_DATA_TEMPR5[53] , \Z\R_DATA_TEMPR5[52] , 
        \Z\R_DATA_TEMPR5[51] , \Z\R_DATA_TEMPR5[50] , 
        \Z\R_DATA_TEMPR5[49] , \Z\R_DATA_TEMPR5[48] , 
        \Z\R_DATA_TEMPR5[47] , \Z\R_DATA_TEMPR5[46] , 
        \Z\R_DATA_TEMPR5[45] , \Z\R_DATA_TEMPR5[44] , 
        \Z\R_DATA_TEMPR5[43] , \Z\R_DATA_TEMPR5[42] , 
        \Z\R_DATA_TEMPR5[41] , \Z\R_DATA_TEMPR5[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[5][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[1] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[1] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_561 (.A(\Z\R_DATA_TEMPR28[29] ), .B(\Z\R_DATA_TEMPR29[29] )
        , .C(\Z\R_DATA_TEMPR30[29] ), .D(\Z\R_DATA_TEMPR31[29] ), .Y(
        OR4_561_Y));
    OR4 OR4_403 (.A(OR4_518_Y), .B(OR2_5_Y), .C(\Z\R_DATA_TEMPR22[40] )
        , .D(\Z\R_DATA_TEMPR23[40] ), .Y(OR4_403_Y));
    OR4 OR4_601 (.A(\Z\R_DATA_TEMPR28[5] ), .B(\Z\R_DATA_TEMPR29[5] ), 
        .C(\Z\R_DATA_TEMPR30[5] ), .D(\Z\R_DATA_TEMPR31[5] ), .Y(
        OR4_601_Y));
    OR2 OR2_68 (.A(\Z\R_DATA_TEMPR20[1] ), .B(\Z\R_DATA_TEMPR21[1] ), 
        .Y(OR2_68_Y));
    OR4 OR4_219 (.A(\Z\R_DATA_TEMPR28[13] ), .B(\Z\R_DATA_TEMPR29[13] )
        , .C(\Z\R_DATA_TEMPR30[13] ), .D(\Z\R_DATA_TEMPR31[13] ), .Y(
        OR4_219_Y));
    OR4 OR4_208 (.A(\Z\R_DATA_TEMPR28[37] ), .B(\Z\R_DATA_TEMPR29[37] )
        , .C(\Z\R_DATA_TEMPR30[37] ), .D(\Z\R_DATA_TEMPR31[37] ), .Y(
        OR4_208_Y));
    OR4 \OR4_R_DATA[68]  (.A(OR4_191_Y), .B(OR4_83_Y), .C(OR4_482_Y), 
        .D(OR4_580_Y), .Y(R_DATA_c[68]));
    OR4 \OR4_R_DATA[19]  (.A(OR4_240_Y), .B(OR4_66_Y), .C(OR4_24_Y), 
        .D(OR4_621_Y), .Y(R_DATA_c[19]));
    OR4 OR4_323 (.A(\Z\R_DATA_TEMPR24[70] ), .B(\Z\R_DATA_TEMPR25[70] )
        , .C(\Z\R_DATA_TEMPR26[70] ), .D(\Z\R_DATA_TEMPR27[70] ), .Y(
        OR4_323_Y));
    OR4 OR4_473 (.A(OR4_370_Y), .B(OR2_23_Y), .C(
        \Z\R_DATA_TEMPR22[77] ), .D(\Z\R_DATA_TEMPR23[77] ), .Y(
        OR4_473_Y));
    OR4 OR4_671 (.A(\Z\R_DATA_TEMPR24[52] ), .B(\Z\R_DATA_TEMPR25[52] )
        , .C(\Z\R_DATA_TEMPR26[52] ), .D(\Z\R_DATA_TEMPR27[52] ), .Y(
        OR4_671_Y));
    OR2 OR2_38 (.A(\Z\R_DATA_TEMPR20[47] ), .B(\Z\R_DATA_TEMPR21[47] ), 
        .Y(OR2_38_Y));
    OR4 \OR4_R_DATA[75]  (.A(OR4_605_Y), .B(OR4_234_Y), .C(OR4_505_Y), 
        .D(OR4_298_Y), .Y(R_DATA_c[75]));
    OR4 OR4_422 (.A(OR4_696_Y), .B(OR4_96_Y), .C(OR4_533_Y), .D(
        OR4_443_Y), .Y(OR4_422_Y));
    OR4 OR4_278 (.A(\Z\R_DATA_TEMPR28[49] ), .B(\Z\R_DATA_TEMPR29[49] )
        , .C(\Z\R_DATA_TEMPR30[49] ), .D(\Z\R_DATA_TEMPR31[49] ), .Y(
        OR4_278_Y));
    OR4 OR4_23 (.A(\Z\R_DATA_TEMPR4[41] ), .B(\Z\R_DATA_TEMPR5[41] ), 
        .C(\Z\R_DATA_TEMPR6[41] ), .D(\Z\R_DATA_TEMPR7[41] ), .Y(
        OR4_23_Y));
    OR4 OR4_199 (.A(\Z\R_DATA_TEMPR0[40] ), .B(\Z\R_DATA_TEMPR1[40] ), 
        .C(\Z\R_DATA_TEMPR2[40] ), .D(\Z\R_DATA_TEMPR3[40] ), .Y(
        OR4_199_Y));
    OR4 OR4_254 (.A(\Z\R_DATA_TEMPR12[3] ), .B(\Z\R_DATA_TEMPR13[3] ), 
        .C(\Z\R_DATA_TEMPR14[3] ), .D(\Z\R_DATA_TEMPR15[3] ), .Y(
        OR4_254_Y));
    OR4 OR4_429 (.A(\Z\R_DATA_TEMPR8[57] ), .B(\Z\R_DATA_TEMPR9[57] ), 
        .C(\Z\R_DATA_TEMPR10[57] ), .D(\Z\R_DATA_TEMPR11[57] ), .Y(
        OR4_429_Y));
    OR4 OR4_262 (.A(\Z\R_DATA_TEMPR0[11] ), .B(\Z\R_DATA_TEMPR1[11] ), 
        .C(\Z\R_DATA_TEMPR2[11] ), .D(\Z\R_DATA_TEMPR3[11] ), .Y(
        OR4_262_Y));
    OR4 OR4_126 (.A(OR4_345_Y), .B(OR2_39_Y), .C(
        \Z\R_DATA_TEMPR22[31] ), .D(\Z\R_DATA_TEMPR23[31] ), .Y(
        OR4_126_Y));
    OR4 OR4_94 (.A(\Z\R_DATA_TEMPR4[65] ), .B(\Z\R_DATA_TEMPR5[65] ), 
        .C(\Z\R_DATA_TEMPR6[65] ), .D(\Z\R_DATA_TEMPR7[65] ), .Y(
        OR4_94_Y));
    OR4 OR4_65 (.A(\Z\R_DATA_TEMPR16[34] ), .B(\Z\R_DATA_TEMPR17[34] ), 
        .C(\Z\R_DATA_TEMPR18[34] ), .D(\Z\R_DATA_TEMPR19[34] ), .Y(
        OR4_65_Y));
    OR4 OR4_360 (.A(\Z\R_DATA_TEMPR16[32] ), .B(\Z\R_DATA_TEMPR17[32] )
        , .C(\Z\R_DATA_TEMPR18[32] ), .D(\Z\R_DATA_TEMPR19[32] ), .Y(
        OR4_360_Y));
    OR4 OR4_355 (.A(\Z\R_DATA_TEMPR16[60] ), .B(\Z\R_DATA_TEMPR17[60] )
        , .C(\Z\R_DATA_TEMPR18[60] ), .D(\Z\R_DATA_TEMPR19[60] ), .Y(
        OR4_355_Y));
    OR4 OR4_344 (.A(\Z\R_DATA_TEMPR28[52] ), .B(\Z\R_DATA_TEMPR29[52] )
        , .C(\Z\R_DATA_TEMPR30[52] ), .D(\Z\R_DATA_TEMPR31[52] ), .Y(
        OR4_344_Y));
    OR4 OR4_328 (.A(\Z\R_DATA_TEMPR8[37] ), .B(\Z\R_DATA_TEMPR9[37] ), 
        .C(\Z\R_DATA_TEMPR10[37] ), .D(\Z\R_DATA_TEMPR11[37] ), .Y(
        OR4_328_Y));
    OR4 OR4_185 (.A(\Z\R_DATA_TEMPR8[43] ), .B(\Z\R_DATA_TEMPR9[43] ), 
        .C(\Z\R_DATA_TEMPR10[43] ), .D(\Z\R_DATA_TEMPR11[43] ), .Y(
        OR4_185_Y));
    OR4 OR4_141 (.A(\Z\R_DATA_TEMPR28[76] ), .B(\Z\R_DATA_TEMPR29[76] )
        , .C(\Z\R_DATA_TEMPR30[76] ), .D(\Z\R_DATA_TEMPR31[76] ), .Y(
        OR4_141_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%25%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0 (
        .A_DOUT({\Z\R_DATA_TEMPR25[39] , \Z\R_DATA_TEMPR25[38] , 
        \Z\R_DATA_TEMPR25[37] , \Z\R_DATA_TEMPR25[36] , 
        \Z\R_DATA_TEMPR25[35] , \Z\R_DATA_TEMPR25[34] , 
        \Z\R_DATA_TEMPR25[33] , \Z\R_DATA_TEMPR25[32] , 
        \Z\R_DATA_TEMPR25[31] , \Z\R_DATA_TEMPR25[30] , 
        \Z\R_DATA_TEMPR25[29] , \Z\R_DATA_TEMPR25[28] , 
        \Z\R_DATA_TEMPR25[27] , \Z\R_DATA_TEMPR25[26] , 
        \Z\R_DATA_TEMPR25[25] , \Z\R_DATA_TEMPR25[24] , 
        \Z\R_DATA_TEMPR25[23] , \Z\R_DATA_TEMPR25[22] , 
        \Z\R_DATA_TEMPR25[21] , \Z\R_DATA_TEMPR25[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR25[19] , \Z\R_DATA_TEMPR25[18] , 
        \Z\R_DATA_TEMPR25[17] , \Z\R_DATA_TEMPR25[16] , 
        \Z\R_DATA_TEMPR25[15] , \Z\R_DATA_TEMPR25[14] , 
        \Z\R_DATA_TEMPR25[13] , \Z\R_DATA_TEMPR25[12] , 
        \Z\R_DATA_TEMPR25[11] , \Z\R_DATA_TEMPR25[10] , 
        \Z\R_DATA_TEMPR25[9] , \Z\R_DATA_TEMPR25[8] , 
        \Z\R_DATA_TEMPR25[7] , \Z\R_DATA_TEMPR25[6] , 
        \Z\R_DATA_TEMPR25[5] , \Z\R_DATA_TEMPR25[4] , 
        \Z\R_DATA_TEMPR25[3] , \Z\R_DATA_TEMPR25[2] , 
        \Z\R_DATA_TEMPR25[1] , \Z\R_DATA_TEMPR25[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[25][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[6] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[6] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[49]  (.A(OR4_607_Y), .B(OR4_440_Y), .C(OR4_395_Y), 
        .D(OR4_278_Y), .Y(R_DATA_c[49]));
    OR4 OR4_717 (.A(\Z\R_DATA_TEMPR28[77] ), .B(\Z\R_DATA_TEMPR29[77] )
        , .C(\Z\R_DATA_TEMPR30[77] ), .D(\Z\R_DATA_TEMPR31[77] ), .Y(
        OR4_717_Y));
    OR4 OR4_36 (.A(\Z\R_DATA_TEMPR8[60] ), .B(\Z\R_DATA_TEMPR9[60] ), 
        .C(\Z\R_DATA_TEMPR10[60] ), .D(\Z\R_DATA_TEMPR11[60] ), .Y(
        OR4_36_Y));
    OR4 OR4_487 (.A(\Z\R_DATA_TEMPR8[76] ), .B(\Z\R_DATA_TEMPR9[76] ), 
        .C(\Z\R_DATA_TEMPR10[76] ), .D(\Z\R_DATA_TEMPR11[76] ), .Y(
        OR4_487_Y));
    OR4 OR4_714 (.A(\Z\R_DATA_TEMPR24[79] ), .B(\Z\R_DATA_TEMPR25[79] )
        , .C(\Z\R_DATA_TEMPR26[79] ), .D(\Z\R_DATA_TEMPR27[79] ), .Y(
        OR4_714_Y));
    OR4 OR4_501 (.A(OR4_397_Y), .B(OR2_47_Y), .C(
        \Z\R_DATA_TEMPR22[17] ), .D(\Z\R_DATA_TEMPR23[17] ), .Y(
        OR4_501_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%27%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0 (
        .A_DOUT({\Z\R_DATA_TEMPR27[39] , \Z\R_DATA_TEMPR27[38] , 
        \Z\R_DATA_TEMPR27[37] , \Z\R_DATA_TEMPR27[36] , 
        \Z\R_DATA_TEMPR27[35] , \Z\R_DATA_TEMPR27[34] , 
        \Z\R_DATA_TEMPR27[33] , \Z\R_DATA_TEMPR27[32] , 
        \Z\R_DATA_TEMPR27[31] , \Z\R_DATA_TEMPR27[30] , 
        \Z\R_DATA_TEMPR27[29] , \Z\R_DATA_TEMPR27[28] , 
        \Z\R_DATA_TEMPR27[27] , \Z\R_DATA_TEMPR27[26] , 
        \Z\R_DATA_TEMPR27[25] , \Z\R_DATA_TEMPR27[24] , 
        \Z\R_DATA_TEMPR27[23] , \Z\R_DATA_TEMPR27[22] , 
        \Z\R_DATA_TEMPR27[21] , \Z\R_DATA_TEMPR27[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR27[19] , \Z\R_DATA_TEMPR27[18] , 
        \Z\R_DATA_TEMPR27[17] , \Z\R_DATA_TEMPR27[16] , 
        \Z\R_DATA_TEMPR27[15] , \Z\R_DATA_TEMPR27[14] , 
        \Z\R_DATA_TEMPR27[13] , \Z\R_DATA_TEMPR27[12] , 
        \Z\R_DATA_TEMPR27[11] , \Z\R_DATA_TEMPR27[10] , 
        \Z\R_DATA_TEMPR27[9] , \Z\R_DATA_TEMPR27[8] , 
        \Z\R_DATA_TEMPR27[7] , \Z\R_DATA_TEMPR27[6] , 
        \Z\R_DATA_TEMPR27[5] , \Z\R_DATA_TEMPR27[4] , 
        \Z\R_DATA_TEMPR27[3] , \Z\R_DATA_TEMPR27[2] , 
        \Z\R_DATA_TEMPR27[1] , \Z\R_DATA_TEMPR27[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[27][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[6] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[6] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_21 (.A(\Z\R_DATA_TEMPR8[63] ), .B(\Z\R_DATA_TEMPR9[63] ), 
        .C(\Z\R_DATA_TEMPR10[63] ), .D(\Z\R_DATA_TEMPR11[63] ), .Y(
        OR4_21_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[3]  (.A(CFG2_5_Y), .B(
        R_ADDR_c[13]), .C(R_EN_c), .Y(\Z\BLKY2[3] ));
    OR4 OR4_129 (.A(\Z\R_DATA_TEMPR24[16] ), .B(\Z\R_DATA_TEMPR25[16] )
        , .C(\Z\R_DATA_TEMPR26[16] ), .D(\Z\R_DATA_TEMPR27[16] ), .Y(
        OR4_129_Y));
    OR4 OR4_571 (.A(OR4_123_Y), .B(OR4_552_Y), .C(OR4_582_Y), .D(
        OR4_237_Y), .Y(OR4_571_Y));
    OR4 OR4_441 (.A(OR4_479_Y), .B(OR2_42_Y), .C(\Z\R_DATA_TEMPR22[8] )
        , .D(\Z\R_DATA_TEMPR23[8] ), .Y(OR4_441_Y));
    OR4 OR4_697 (.A(\Z\R_DATA_TEMPR28[61] ), .B(\Z\R_DATA_TEMPR29[61] )
        , .C(\Z\R_DATA_TEMPR30[61] ), .D(\Z\R_DATA_TEMPR31[61] ), .Y(
        OR4_697_Y));
    OR4 OR4_448 (.A(\Z\R_DATA_TEMPR28[42] ), .B(\Z\R_DATA_TEMPR29[42] )
        , .C(\Z\R_DATA_TEMPR30[42] ), .D(\Z\R_DATA_TEMPR31[42] ), .Y(
        OR4_448_Y));
    OR4 OR4_285 (.A(\Z\R_DATA_TEMPR16[33] ), .B(\Z\R_DATA_TEMPR17[33] )
        , .C(\Z\R_DATA_TEMPR18[33] ), .D(\Z\R_DATA_TEMPR19[33] ), .Y(
        OR4_285_Y));
    OR4 OR4_202 (.A(\Z\R_DATA_TEMPR24[39] ), .B(\Z\R_DATA_TEMPR25[39] )
        , .C(\Z\R_DATA_TEMPR26[39] ), .D(\Z\R_DATA_TEMPR27[39] ), .Y(
        OR4_202_Y));
    OR4 \OR4_R_DATA[69]  (.A(OR4_439_Y), .B(OR4_286_Y), .C(OR4_253_Y), 
        .D(OR4_103_Y), .Y(R_DATA_c[69]));
    OR4 OR4_655 (.A(\Z\R_DATA_TEMPR16[59] ), .B(\Z\R_DATA_TEMPR17[59] )
        , .C(\Z\R_DATA_TEMPR18[59] ), .D(\Z\R_DATA_TEMPR19[59] ), .Y(
        OR4_655_Y));
    OR4 OR4_272 (.A(\Z\R_DATA_TEMPR24[18] ), .B(\Z\R_DATA_TEMPR25[18] )
        , .C(\Z\R_DATA_TEMPR26[18] ), .D(\Z\R_DATA_TEMPR27[18] ), .Y(
        OR4_272_Y));
    OR4 OR4_565 (.A(\Z\R_DATA_TEMPR0[45] ), .B(\Z\R_DATA_TEMPR1[45] ), 
        .C(\Z\R_DATA_TEMPR2[45] ), .D(\Z\R_DATA_TEMPR3[45] ), .Y(
        OR4_565_Y));
    OR4 OR4_44 (.A(OR4_461_Y), .B(OR2_2_Y), .C(\Z\R_DATA_TEMPR22[52] ), 
        .D(\Z\R_DATA_TEMPR23[52] ), .Y(OR4_44_Y));
    OR4 OR4_549 (.A(\Z\R_DATA_TEMPR4[30] ), .B(\Z\R_DATA_TEMPR5[30] ), 
        .C(\Z\R_DATA_TEMPR6[30] ), .D(\Z\R_DATA_TEMPR7[30] ), .Y(
        OR4_549_Y));
    OR4 OR4_435 (.A(\Z\R_DATA_TEMPR24[63] ), .B(\Z\R_DATA_TEMPR25[63] )
        , .C(\Z\R_DATA_TEMPR26[63] ), .D(\Z\R_DATA_TEMPR27[63] ), .Y(
        OR4_435_Y));
    OR4 OR4_300 (.A(OR4_406_Y), .B(OR2_11_Y), .C(
        \Z\R_DATA_TEMPR22[50] ), .D(\Z\R_DATA_TEMPR23[50] ), .Y(
        OR4_300_Y));
    OR4 OR4_540 (.A(\Z\R_DATA_TEMPR4[31] ), .B(\Z\R_DATA_TEMPR5[31] ), 
        .C(\Z\R_DATA_TEMPR6[31] ), .D(\Z\R_DATA_TEMPR7[31] ), .Y(
        OR4_540_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[0]  (.A(CFG2_4_Y), .B(
        W_ADDR_c[13]), .C(W_EN_c), .Y(\Z\BLKX2[0] ));
    OR4 OR4_483 (.A(\Z\R_DATA_TEMPR16[58] ), .B(\Z\R_DATA_TEMPR17[58] )
        , .C(\Z\R_DATA_TEMPR18[58] ), .D(\Z\R_DATA_TEMPR19[58] ), .Y(
        OR4_483_Y));
    OR4 OR4_681 (.A(\Z\R_DATA_TEMPR24[29] ), .B(\Z\R_DATA_TEMPR25[29] )
        , .C(\Z\R_DATA_TEMPR26[29] ), .D(\Z\R_DATA_TEMPR27[29] ), .Y(
        OR4_681_Y));
    OR4 OR4_663 (.A(\Z\R_DATA_TEMPR12[45] ), .B(\Z\R_DATA_TEMPR13[45] )
        , .C(\Z\R_DATA_TEMPR14[45] ), .D(\Z\R_DATA_TEMPR15[45] ), .Y(
        OR4_663_Y));
    OR4 OR4_370 (.A(\Z\R_DATA_TEMPR16[77] ), .B(\Z\R_DATA_TEMPR17[77] )
        , .C(\Z\R_DATA_TEMPR18[77] ), .D(\Z\R_DATA_TEMPR19[77] ), .Y(
        OR4_370_Y));
    OR4 OR4_288 (.A(\Z\R_DATA_TEMPR8[29] ), .B(\Z\R_DATA_TEMPR9[29] ), 
        .C(\Z\R_DATA_TEMPR10[29] ), .D(\Z\R_DATA_TEMPR11[29] ), .Y(
        OR4_288_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%29%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C1 (
        .A_DOUT({\Z\R_DATA_TEMPR29[79] , \Z\R_DATA_TEMPR29[78] , 
        \Z\R_DATA_TEMPR29[77] , \Z\R_DATA_TEMPR29[76] , 
        \Z\R_DATA_TEMPR29[75] , \Z\R_DATA_TEMPR29[74] , 
        \Z\R_DATA_TEMPR29[73] , \Z\R_DATA_TEMPR29[72] , 
        \Z\R_DATA_TEMPR29[71] , \Z\R_DATA_TEMPR29[70] , 
        \Z\R_DATA_TEMPR29[69] , \Z\R_DATA_TEMPR29[68] , 
        \Z\R_DATA_TEMPR29[67] , \Z\R_DATA_TEMPR29[66] , 
        \Z\R_DATA_TEMPR29[65] , \Z\R_DATA_TEMPR29[64] , 
        \Z\R_DATA_TEMPR29[63] , \Z\R_DATA_TEMPR29[62] , 
        \Z\R_DATA_TEMPR29[61] , \Z\R_DATA_TEMPR29[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR29[59] , \Z\R_DATA_TEMPR29[58] , 
        \Z\R_DATA_TEMPR29[57] , \Z\R_DATA_TEMPR29[56] , 
        \Z\R_DATA_TEMPR29[55] , \Z\R_DATA_TEMPR29[54] , 
        \Z\R_DATA_TEMPR29[53] , \Z\R_DATA_TEMPR29[52] , 
        \Z\R_DATA_TEMPR29[51] , \Z\R_DATA_TEMPR29[50] , 
        \Z\R_DATA_TEMPR29[49] , \Z\R_DATA_TEMPR29[48] , 
        \Z\R_DATA_TEMPR29[47] , \Z\R_DATA_TEMPR29[46] , 
        \Z\R_DATA_TEMPR29[45] , \Z\R_DATA_TEMPR29[44] , 
        \Z\R_DATA_TEMPR29[43] , \Z\R_DATA_TEMPR29[42] , 
        \Z\R_DATA_TEMPR29[41] , \Z\R_DATA_TEMPR29[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[29][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[7] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[7] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[54]  (.A(OR4_247_Y), .B(OR4_708_Y), .C(OR4_324_Y), 
        .D(OR4_650_Y), .Y(R_DATA_c[54]));
    OR4 OR4_30 (.A(\Z\R_DATA_TEMPR0[60] ), .B(\Z\R_DATA_TEMPR1[60] ), 
        .C(\Z\R_DATA_TEMPR2[60] ), .D(\Z\R_DATA_TEMPR3[60] ), .Y(
        OR4_30_Y));
    OR4 OR4_650 (.A(\Z\R_DATA_TEMPR28[54] ), .B(\Z\R_DATA_TEMPR29[54] )
        , .C(\Z\R_DATA_TEMPR30[54] ), .D(\Z\R_DATA_TEMPR31[54] ), .Y(
        OR4_650_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%9%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C1 (
        .A_DOUT({\Z\R_DATA_TEMPR9[79] , \Z\R_DATA_TEMPR9[78] , 
        \Z\R_DATA_TEMPR9[77] , \Z\R_DATA_TEMPR9[76] , 
        \Z\R_DATA_TEMPR9[75] , \Z\R_DATA_TEMPR9[74] , 
        \Z\R_DATA_TEMPR9[73] , \Z\R_DATA_TEMPR9[72] , 
        \Z\R_DATA_TEMPR9[71] , \Z\R_DATA_TEMPR9[70] , 
        \Z\R_DATA_TEMPR9[69] , \Z\R_DATA_TEMPR9[68] , 
        \Z\R_DATA_TEMPR9[67] , \Z\R_DATA_TEMPR9[66] , 
        \Z\R_DATA_TEMPR9[65] , \Z\R_DATA_TEMPR9[64] , 
        \Z\R_DATA_TEMPR9[63] , \Z\R_DATA_TEMPR9[62] , 
        \Z\R_DATA_TEMPR9[61] , \Z\R_DATA_TEMPR9[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR9[59] , \Z\R_DATA_TEMPR9[58] , 
        \Z\R_DATA_TEMPR9[57] , \Z\R_DATA_TEMPR9[56] , 
        \Z\R_DATA_TEMPR9[55] , \Z\R_DATA_TEMPR9[54] , 
        \Z\R_DATA_TEMPR9[53] , \Z\R_DATA_TEMPR9[52] , 
        \Z\R_DATA_TEMPR9[51] , \Z\R_DATA_TEMPR9[50] , 
        \Z\R_DATA_TEMPR9[49] , \Z\R_DATA_TEMPR9[48] , 
        \Z\R_DATA_TEMPR9[47] , \Z\R_DATA_TEMPR9[46] , 
        \Z\R_DATA_TEMPR9[45] , \Z\R_DATA_TEMPR9[44] , 
        \Z\R_DATA_TEMPR9[43] , \Z\R_DATA_TEMPR9[42] , 
        \Z\R_DATA_TEMPR9[41] , \Z\R_DATA_TEMPR9[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[9][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[2] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[2] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_627 (.A(OR4_343_Y), .B(OR2_8_Y), .C(\Z\R_DATA_TEMPR22[45] )
        , .D(\Z\R_DATA_TEMPR23[45] ), .Y(OR4_627_Y));
    OR4 OR4_297 (.A(\Z\R_DATA_TEMPR4[22] ), .B(\Z\R_DATA_TEMPR5[22] ), 
        .C(\Z\R_DATA_TEMPR6[22] ), .D(\Z\R_DATA_TEMPR7[22] ), .Y(
        OR4_297_Y));
    OR4 OR4_37 (.A(OR4_703_Y), .B(OR4_549_Y), .C(OR4_711_Y), .D(
        OR4_311_Y), .Y(OR4_37_Y));
    OR4 OR4_197 (.A(\Z\R_DATA_TEMPR12[23] ), .B(\Z\R_DATA_TEMPR13[23] )
        , .C(\Z\R_DATA_TEMPR14[23] ), .D(\Z\R_DATA_TEMPR15[23] ), .Y(
        OR4_197_Y));
    OR4 OR4_357 (.A(\Z\R_DATA_TEMPR16[79] ), .B(\Z\R_DATA_TEMPR17[79] )
        , .C(\Z\R_DATA_TEMPR18[79] ), .D(\Z\R_DATA_TEMPR19[79] ), .Y(
        OR4_357_Y));
    OR4 OR4_150 (.A(\Z\R_DATA_TEMPR16[71] ), .B(\Z\R_DATA_TEMPR17[71] )
        , .C(\Z\R_DATA_TEMPR18[71] ), .D(\Z\R_DATA_TEMPR19[71] ), .Y(
        OR4_150_Y));
    OR4 OR4_434 (.A(OR4_679_Y), .B(OR4_541_Y), .C(OR4_528_Y), .D(
        OR4_260_Y), .Y(OR4_434_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[5]  (.A(CFG2_6_Y), .B(
        R_ADDR_c[13]), .C(R_EN_c), .Y(\Z\BLKY2[5] ));
    CFG2 #( .INIT(4'h2) )  CFG2_7 (.A(W_ADDR_c[12]), .B(W_ADDR_c[11]), 
        .Y(CFG2_7_Y));
    OR4 OR4_163 (.A(\Z\R_DATA_TEMPR28[59] ), .B(\Z\R_DATA_TEMPR29[59] )
        , .C(\Z\R_DATA_TEMPR30[59] ), .D(\Z\R_DATA_TEMPR31[59] ), .Y(
        OR4_163_Y));
    OR4 OR4_343 (.A(\Z\R_DATA_TEMPR16[45] ), .B(\Z\R_DATA_TEMPR17[45] )
        , .C(\Z\R_DATA_TEMPR18[45] ), .D(\Z\R_DATA_TEMPR19[45] ), .Y(
        OR4_343_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[7]  (.A(CFG2_5_Y), .B(
        R_ADDR_c[13]), .C(R_EN_c), .Y(\Z\BLKY2[7] ));
    OR4 OR4_336 (.A(OR4_655_Y), .B(OR2_54_Y), .C(
        \Z\R_DATA_TEMPR22[59] ), .D(\Z\R_DATA_TEMPR23[59] ), .Y(
        OR4_336_Y));
    OR4 OR4_415 (.A(\Z\R_DATA_TEMPR0[31] ), .B(\Z\R_DATA_TEMPR1[31] ), 
        .C(\Z\R_DATA_TEMPR2[31] ), .D(\Z\R_DATA_TEMPR3[31] ), .Y(
        OR4_415_Y));
    OR4 OR4_442 (.A(\Z\R_DATA_TEMPR16[51] ), .B(\Z\R_DATA_TEMPR17[51] )
        , .C(\Z\R_DATA_TEMPR18[51] ), .D(\Z\R_DATA_TEMPR19[51] ), .Y(
        OR4_442_Y));
    OR4 OR4_294 (.A(\Z\R_DATA_TEMPR28[57] ), .B(\Z\R_DATA_TEMPR29[57] )
        , .C(\Z\R_DATA_TEMPR30[57] ), .D(\Z\R_DATA_TEMPR31[57] ), .Y(
        OR4_294_Y));
    OR4 OR4_449 (.A(\Z\R_DATA_TEMPR12[35] ), .B(\Z\R_DATA_TEMPR13[35] )
        , .C(\Z\R_DATA_TEMPR14[35] ), .D(\Z\R_DATA_TEMPR15[35] ), .Y(
        OR4_449_Y));
    OR4 OR4_505 (.A(\Z\R_DATA_TEMPR24[75] ), .B(\Z\R_DATA_TEMPR25[75] )
        , .C(\Z\R_DATA_TEMPR26[75] ), .D(\Z\R_DATA_TEMPR27[75] ), .Y(
        OR4_505_Y));
    OR4 \OR4_R_DATA[24]  (.A(OR4_630_Y), .B(OR4_374_Y), .C(OR4_4_Y), 
        .D(OR4_315_Y), .Y(R_DATA_c[24]));
    OR4 OR4_85 (.A(\Z\R_DATA_TEMPR12[39] ), .B(\Z\R_DATA_TEMPR13[39] ), 
        .C(\Z\R_DATA_TEMPR14[39] ), .D(\Z\R_DATA_TEMPR15[39] ), .Y(
        OR4_85_Y));
    OR4 \OR4_R_DATA[12]  (.A(OR4_526_Y), .B(OR4_502_Y), .C(OR4_398_Y), 
        .D(OR4_69_Y), .Y(R_DATA_c[12]));
    OR4 OR4_158 (.A(\Z\R_DATA_TEMPR4[57] ), .B(\Z\R_DATA_TEMPR5[57] ), 
        .C(\Z\R_DATA_TEMPR6[57] ), .D(\Z\R_DATA_TEMPR7[57] ), .Y(
        OR4_158_Y));
    OR4 OR4_146 (.A(\Z\R_DATA_TEMPR16[76] ), .B(\Z\R_DATA_TEMPR17[76] )
        , .C(\Z\R_DATA_TEMPR18[76] ), .D(\Z\R_DATA_TEMPR19[76] ), .Y(
        OR4_146_Y));
    OR4 \OR4_R_DATA[78]  (.A(OR4_662_Y), .B(OR4_564_Y), .C(OR4_248_Y), 
        .D(OR4_326_Y), .Y(R_DATA_c[78]));
    OR4 OR4_581 (.A(\Z\R_DATA_TEMPR12[74] ), .B(\Z\R_DATA_TEMPR13[74] )
        , .C(\Z\R_DATA_TEMPR14[74] ), .D(\Z\R_DATA_TEMPR15[74] ), .Y(
        OR4_581_Y));
    OR4 OR4_575 (.A(\Z\R_DATA_TEMPR4[5] ), .B(\Z\R_DATA_TEMPR5[5] ), 
        .C(\Z\R_DATA_TEMPR6[5] ), .D(\Z\R_DATA_TEMPR7[5] ), .Y(
        OR4_575_Y));
    OR2 OR2_45 (.A(\Z\R_DATA_TEMPR20[57] ), .B(\Z\R_DATA_TEMPR21[57] ), 
        .Y(OR2_45_Y));
    OR4 OR4_69 (.A(\Z\R_DATA_TEMPR28[12] ), .B(\Z\R_DATA_TEMPR29[12] ), 
        .C(\Z\R_DATA_TEMPR30[12] ), .D(\Z\R_DATA_TEMPR31[12] ), .Y(
        OR4_69_Y));
    OR4 OR4_603 (.A(\Z\R_DATA_TEMPR24[43] ), .B(\Z\R_DATA_TEMPR25[43] )
        , .C(\Z\R_DATA_TEMPR26[43] ), .D(\Z\R_DATA_TEMPR27[43] ), .Y(
        OR4_603_Y));
    OR2 OR2_56 (.A(\Z\R_DATA_TEMPR20[21] ), .B(\Z\R_DATA_TEMPR21[21] ), 
        .Y(OR2_56_Y));
    OR4 OR4_227 (.A(\Z\R_DATA_TEMPR12[73] ), .B(\Z\R_DATA_TEMPR13[73] )
        , .C(\Z\R_DATA_TEMPR14[73] ), .D(\Z\R_DATA_TEMPR15[73] ), .Y(
        OR4_227_Y));
    OR4 OR4_673 (.A(OR4_104_Y), .B(OR2_9_Y), .C(\Z\R_DATA_TEMPR22[26] )
        , .D(\Z\R_DATA_TEMPR23[26] ), .Y(OR4_673_Y));
    OR4 OR4_395 (.A(\Z\R_DATA_TEMPR24[49] ), .B(\Z\R_DATA_TEMPR25[49] )
        , .C(\Z\R_DATA_TEMPR26[49] ), .D(\Z\R_DATA_TEMPR27[49] ), .Y(
        OR4_395_Y));
    OR4 OR4_414 (.A(\Z\R_DATA_TEMPR12[50] ), .B(\Z\R_DATA_TEMPR13[50] )
        , .C(\Z\R_DATA_TEMPR14[50] ), .D(\Z\R_DATA_TEMPR15[50] ), .Y(
        OR4_414_Y));
    OR4 OR4_127 (.A(\Z\R_DATA_TEMPR8[65] ), .B(\Z\R_DATA_TEMPR9[65] ), 
        .C(\Z\R_DATA_TEMPR10[65] ), .D(\Z\R_DATA_TEMPR11[65] ), .Y(
        OR4_127_Y));
    OR4 OR4_348 (.A(\Z\R_DATA_TEMPR28[74] ), .B(\Z\R_DATA_TEMPR29[74] )
        , .C(\Z\R_DATA_TEMPR30[74] ), .D(\Z\R_DATA_TEMPR31[74] ), .Y(
        OR4_348_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%30%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C1 (
        .A_DOUT({\Z\R_DATA_TEMPR30[79] , \Z\R_DATA_TEMPR30[78] , 
        \Z\R_DATA_TEMPR30[77] , \Z\R_DATA_TEMPR30[76] , 
        \Z\R_DATA_TEMPR30[75] , \Z\R_DATA_TEMPR30[74] , 
        \Z\R_DATA_TEMPR30[73] , \Z\R_DATA_TEMPR30[72] , 
        \Z\R_DATA_TEMPR30[71] , \Z\R_DATA_TEMPR30[70] , 
        \Z\R_DATA_TEMPR30[69] , \Z\R_DATA_TEMPR30[68] , 
        \Z\R_DATA_TEMPR30[67] , \Z\R_DATA_TEMPR30[66] , 
        \Z\R_DATA_TEMPR30[65] , \Z\R_DATA_TEMPR30[64] , 
        \Z\R_DATA_TEMPR30[63] , \Z\R_DATA_TEMPR30[62] , 
        \Z\R_DATA_TEMPR30[61] , \Z\R_DATA_TEMPR30[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR30[59] , \Z\R_DATA_TEMPR30[58] , 
        \Z\R_DATA_TEMPR30[57] , \Z\R_DATA_TEMPR30[56] , 
        \Z\R_DATA_TEMPR30[55] , \Z\R_DATA_TEMPR30[54] , 
        \Z\R_DATA_TEMPR30[53] , \Z\R_DATA_TEMPR30[52] , 
        \Z\R_DATA_TEMPR30[51] , \Z\R_DATA_TEMPR30[50] , 
        \Z\R_DATA_TEMPR30[49] , \Z\R_DATA_TEMPR30[48] , 
        \Z\R_DATA_TEMPR30[47] , \Z\R_DATA_TEMPR30[46] , 
        \Z\R_DATA_TEMPR30[45] , \Z\R_DATA_TEMPR30[44] , 
        \Z\R_DATA_TEMPR30[43] , \Z\R_DATA_TEMPR30[42] , 
        \Z\R_DATA_TEMPR30[41] , \Z\R_DATA_TEMPR30[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[30][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[7] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[7] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_162 (.A(\Z\R_DATA_TEMPR12[47] ), .B(\Z\R_DATA_TEMPR13[47] )
        , .C(\Z\R_DATA_TEMPR14[47] ), .D(\Z\R_DATA_TEMPR15[47] ), .Y(
        OR4_162_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%16%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0 (
        .A_DOUT({\Z\R_DATA_TEMPR16[39] , \Z\R_DATA_TEMPR16[38] , 
        \Z\R_DATA_TEMPR16[37] , \Z\R_DATA_TEMPR16[36] , 
        \Z\R_DATA_TEMPR16[35] , \Z\R_DATA_TEMPR16[34] , 
        \Z\R_DATA_TEMPR16[33] , \Z\R_DATA_TEMPR16[32] , 
        \Z\R_DATA_TEMPR16[31] , \Z\R_DATA_TEMPR16[30] , 
        \Z\R_DATA_TEMPR16[29] , \Z\R_DATA_TEMPR16[28] , 
        \Z\R_DATA_TEMPR16[27] , \Z\R_DATA_TEMPR16[26] , 
        \Z\R_DATA_TEMPR16[25] , \Z\R_DATA_TEMPR16[24] , 
        \Z\R_DATA_TEMPR16[23] , \Z\R_DATA_TEMPR16[22] , 
        \Z\R_DATA_TEMPR16[21] , \Z\R_DATA_TEMPR16[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR16[19] , \Z\R_DATA_TEMPR16[18] , 
        \Z\R_DATA_TEMPR16[17] , \Z\R_DATA_TEMPR16[16] , 
        \Z\R_DATA_TEMPR16[15] , \Z\R_DATA_TEMPR16[14] , 
        \Z\R_DATA_TEMPR16[13] , \Z\R_DATA_TEMPR16[12] , 
        \Z\R_DATA_TEMPR16[11] , \Z\R_DATA_TEMPR16[10] , 
        \Z\R_DATA_TEMPR16[9] , \Z\R_DATA_TEMPR16[8] , 
        \Z\R_DATA_TEMPR16[7] , \Z\R_DATA_TEMPR16[6] , 
        \Z\R_DATA_TEMPR16[5] , \Z\R_DATA_TEMPR16[4] , 
        \Z\R_DATA_TEMPR16[3] , \Z\R_DATA_TEMPR16[2] , 
        \Z\R_DATA_TEMPR16[1] , \Z\R_DATA_TEMPR16[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[16][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[4] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[4] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_282 (.A(OR4_565_Y), .B(OR4_271_Y), .C(OR4_291_Y), .D(
        OR4_663_Y), .Y(OR4_282_Y));
    OR4 OR4_316 (.A(OR4_379_Y), .B(OR4_53_Y), .C(OR4_328_Y), .D(
        OR4_678_Y), .Y(OR4_316_Y));
    OR2 OR2_65 (.A(\Z\R_DATA_TEMPR20[39] ), .B(\Z\R_DATA_TEMPR21[39] ), 
        .Y(OR2_65_Y));
    OR4 OR4_134 (.A(\Z\R_DATA_TEMPR12[69] ), .B(\Z\R_DATA_TEMPR13[69] )
        , .C(\Z\R_DATA_TEMPR14[69] ), .D(\Z\R_DATA_TEMPR15[69] ), .Y(
        OR4_134_Y));
    OR2 OR2_35 (.A(\Z\R_DATA_TEMPR20[22] ), .B(\Z\R_DATA_TEMPR21[22] ), 
        .Y(OR2_35_Y));
    OR4 OR4_103 (.A(\Z\R_DATA_TEMPR28[69] ), .B(\Z\R_DATA_TEMPR29[69] )
        , .C(\Z\R_DATA_TEMPR30[69] ), .D(\Z\R_DATA_TEMPR31[69] ), .Y(
        OR4_103_Y));
    OR4 OR4_224 (.A(\Z\R_DATA_TEMPR0[3] ), .B(\Z\R_DATA_TEMPR1[3] ), 
        .C(\Z\R_DATA_TEMPR2[3] ), .D(\Z\R_DATA_TEMPR3[3] ), .Y(
        OR4_224_Y));
    OR4 OR4_149 (.A(\Z\R_DATA_TEMPR4[8] ), .B(\Z\R_DATA_TEMPR5[8] ), 
        .C(\Z\R_DATA_TEMPR6[8] ), .D(\Z\R_DATA_TEMPR7[8] ), .Y(
        OR4_149_Y));
    OR4 OR4_380 (.A(\Z\R_DATA_TEMPR28[14] ), .B(\Z\R_DATA_TEMPR29[14] )
        , .C(\Z\R_DATA_TEMPR30[14] ), .D(\Z\R_DATA_TEMPR31[14] ), .Y(
        OR4_380_Y));
    OR4 \OR4_R_DATA[13]  (.A(OR4_434_Y), .B(OR4_266_Y), .C(OR4_236_Y), 
        .D(OR4_219_Y), .Y(R_DATA_c[13]));
    OR4 OR4_173 (.A(\Z\R_DATA_TEMPR28[16] ), .B(\Z\R_DATA_TEMPR29[16] )
        , .C(\Z\R_DATA_TEMPR30[16] ), .D(\Z\R_DATA_TEMPR31[16] ), .Y(
        OR4_173_Y));
    OR4 \OR4_R_DATA[42]  (.A(OR4_183_Y), .B(OR4_156_Y), .C(OR4_49_Y), 
        .D(OR4_448_Y), .Y(R_DATA_c[42]));
    OR4 OR4_269 (.A(\Z\R_DATA_TEMPR12[75] ), .B(\Z\R_DATA_TEMPR13[75] )
        , .C(\Z\R_DATA_TEMPR14[75] ), .D(\Z\R_DATA_TEMPR15[75] ), .Y(
        OR4_269_Y));
    OR4 OR4_695 (.A(\Z\R_DATA_TEMPR16[15] ), .B(\Z\R_DATA_TEMPR17[15] )
        , .C(\Z\R_DATA_TEMPR18[15] ), .D(\Z\R_DATA_TEMPR19[15] ), .Y(
        OR4_695_Y));
    OR4 OR4_62 (.A(OR4_216_Y), .B(OR4_625_Y), .C(OR4_51_Y), .D(
        OR4_411_Y), .Y(OR4_62_Y));
    OR4 OR4_38 (.A(OR4_377_Y), .B(OR2_37_Y), .C(\Z\R_DATA_TEMPR22[38] )
        , .D(\Z\R_DATA_TEMPR23[38] ), .Y(OR4_38_Y));
    OR4 OR4_325 (.A(\Z\R_DATA_TEMPR0[43] ), .B(\Z\R_DATA_TEMPR1[43] ), 
        .C(\Z\R_DATA_TEMPR2[43] ), .D(\Z\R_DATA_TEMPR3[43] ), .Y(
        OR4_325_Y));
    OR4 OR4_536 (.A(OR4_148_Y), .B(OR2_52_Y), .C(
        \Z\R_DATA_TEMPR22[28] ), .D(\Z\R_DATA_TEMPR23[28] ), .Y(
        OR4_536_Y));
    OR2 OR2_50 (.A(\Z\R_DATA_TEMPR20[60] ), .B(\Z\R_DATA_TEMPR21[60] ), 
        .Y(OR2_50_Y));
    OR4 \OR4_R_DATA[62]  (.A(OR4_19_Y), .B(OR4_716_Y), .C(OR4_618_Y), 
        .D(OR4_292_Y), .Y(R_DATA_c[62]));
    OR4 OR4_114 (.A(\Z\R_DATA_TEMPR4[46] ), .B(\Z\R_DATA_TEMPR5[46] ), 
        .C(\Z\R_DATA_TEMPR6[46] ), .D(\Z\R_DATA_TEMPR7[46] ), .Y(
        OR4_114_Y));
    OR4 OR4_155 (.A(\Z\R_DATA_TEMPR4[55] ), .B(\Z\R_DATA_TEMPR5[55] ), 
        .C(\Z\R_DATA_TEMPR6[55] ), .D(\Z\R_DATA_TEMPR7[55] ), .Y(
        OR4_155_Y));
    OR4 \OR4_R_DATA[79]  (.A(OR4_218_Y), .B(OR4_42_Y), .C(OR4_714_Y), 
        .D(OR4_595_Y), .Y(R_DATA_c[79]));
    OR2 OR2_57 (.A(\Z\R_DATA_TEMPR20[73] ), .B(\Z\R_DATA_TEMPR21[73] ), 
        .Y(OR2_57_Y));
    OR4 OR4_457 (.A(\Z\R_DATA_TEMPR24[5] ), .B(\Z\R_DATA_TEMPR25[5] ), 
        .C(\Z\R_DATA_TEMPR26[5] ), .D(\Z\R_DATA_TEMPR27[5] ), .Y(
        OR4_457_Y));
    OR4 OR4_102 (.A(\Z\R_DATA_TEMPR16[70] ), .B(\Z\R_DATA_TEMPR17[70] )
        , .C(\Z\R_DATA_TEMPR18[70] ), .D(\Z\R_DATA_TEMPR19[70] ), .Y(
        OR4_102_Y));
    INV \INVBLKY0[0]  (.A(R_ADDR_c[9]), .Y(\Z\BLKY0[0] ));
    OR4 OR4_690 (.A(OR4_91_Y), .B(OR4_527_Y), .C(OR4_675_Y), .D(
        OR4_310_Y), .Y(OR4_690_Y));
    OR4 OR4_172 (.A(\Z\R_DATA_TEMPR12[28] ), .B(\Z\R_DATA_TEMPR13[28] )
        , .C(\Z\R_DATA_TEMPR14[28] ), .D(\Z\R_DATA_TEMPR15[28] ), .Y(
        OR4_172_Y));
    OR4 \OR4_R_DATA[51]  (.A(OR4_277_Y), .B(OR4_250_Y), .C(OR4_261_Y), 
        .D(OR4_25_Y), .Y(R_DATA_c[51]));
    OR4 \OR4_R_DATA[43]  (.A(OR4_88_Y), .B(OR4_628_Y), .C(OR4_603_Y), 
        .D(OR4_577_Y), .Y(R_DATA_c[43]));
    OR4 OR4_647 (.A(\Z\R_DATA_TEMPR24[21] ), .B(\Z\R_DATA_TEMPR25[21] )
        , .C(\Z\R_DATA_TEMPR26[21] ), .D(\Z\R_DATA_TEMPR27[21] ), .Y(
        OR4_647_Y));
    OR4 OR4_711 (.A(\Z\R_DATA_TEMPR8[30] ), .B(\Z\R_DATA_TEMPR9[30] ), 
        .C(\Z\R_DATA_TEMPR10[30] ), .D(\Z\R_DATA_TEMPR11[30] ), .Y(
        OR4_711_Y));
    OR4 OR4_585 (.A(\Z\R_DATA_TEMPR12[29] ), .B(\Z\R_DATA_TEMPR13[29] )
        , .C(\Z\R_DATA_TEMPR14[29] ), .D(\Z\R_DATA_TEMPR15[29] ), .Y(
        OR4_585_Y));
    OR4 OR4_255 (.A(\Z\R_DATA_TEMPR28[32] ), .B(\Z\R_DATA_TEMPR29[32] )
        , .C(\Z\R_DATA_TEMPR30[32] ), .D(\Z\R_DATA_TEMPR31[32] ), .Y(
        OR4_255_Y));
    OR4 OR4_397 (.A(\Z\R_DATA_TEMPR16[17] ), .B(\Z\R_DATA_TEMPR17[17] )
        , .C(\Z\R_DATA_TEMPR18[17] ), .D(\Z\R_DATA_TEMPR19[17] ), .Y(
        OR4_397_Y));
    OR4 OR4_190 (.A(\Z\R_DATA_TEMPR16[78] ), .B(\Z\R_DATA_TEMPR17[78] )
        , .C(\Z\R_DATA_TEMPR18[78] ), .D(\Z\R_DATA_TEMPR19[78] ), .Y(
        OR4_190_Y));
    OR4 OR4_625 (.A(\Z\R_DATA_TEMPR4[52] ), .B(\Z\R_DATA_TEMPR5[52] ), 
        .C(\Z\R_DATA_TEMPR6[52] ), .D(\Z\R_DATA_TEMPR7[52] ), .Y(
        OR4_625_Y));
    OR4 OR4_538 (.A(\Z\R_DATA_TEMPR8[31] ), .B(\Z\R_DATA_TEMPR9[31] ), 
        .C(\Z\R_DATA_TEMPR10[31] ), .D(\Z\R_DATA_TEMPR11[31] ), .Y(
        OR4_538_Y));
    OR4 OR4_26 (.A(\Z\R_DATA_TEMPR28[20] ), .B(\Z\R_DATA_TEMPR29[20] ), 
        .C(\Z\R_DATA_TEMPR30[20] ), .D(\Z\R_DATA_TEMPR31[20] ), .Y(
        OR4_26_Y));
    OR4 OR4_53 (.A(\Z\R_DATA_TEMPR4[37] ), .B(\Z\R_DATA_TEMPR5[37] ), 
        .C(\Z\R_DATA_TEMPR6[37] ), .D(\Z\R_DATA_TEMPR7[37] ), .Y(
        OR4_53_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%0%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C1 (
        .A_DOUT({\Z\R_DATA_TEMPR0[79] , \Z\R_DATA_TEMPR0[78] , 
        \Z\R_DATA_TEMPR0[77] , \Z\R_DATA_TEMPR0[76] , 
        \Z\R_DATA_TEMPR0[75] , \Z\R_DATA_TEMPR0[74] , 
        \Z\R_DATA_TEMPR0[73] , \Z\R_DATA_TEMPR0[72] , 
        \Z\R_DATA_TEMPR0[71] , \Z\R_DATA_TEMPR0[70] , 
        \Z\R_DATA_TEMPR0[69] , \Z\R_DATA_TEMPR0[68] , 
        \Z\R_DATA_TEMPR0[67] , \Z\R_DATA_TEMPR0[66] , 
        \Z\R_DATA_TEMPR0[65] , \Z\R_DATA_TEMPR0[64] , 
        \Z\R_DATA_TEMPR0[63] , \Z\R_DATA_TEMPR0[62] , 
        \Z\R_DATA_TEMPR0[61] , \Z\R_DATA_TEMPR0[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR0[59] , \Z\R_DATA_TEMPR0[58] , 
        \Z\R_DATA_TEMPR0[57] , \Z\R_DATA_TEMPR0[56] , 
        \Z\R_DATA_TEMPR0[55] , \Z\R_DATA_TEMPR0[54] , 
        \Z\R_DATA_TEMPR0[53] , \Z\R_DATA_TEMPR0[52] , 
        \Z\R_DATA_TEMPR0[51] , \Z\R_DATA_TEMPR0[50] , 
        \Z\R_DATA_TEMPR0[49] , \Z\R_DATA_TEMPR0[48] , 
        \Z\R_DATA_TEMPR0[47] , \Z\R_DATA_TEMPR0[46] , 
        \Z\R_DATA_TEMPR0[45] , \Z\R_DATA_TEMPR0[44] , 
        \Z\R_DATA_TEMPR0[43] , \Z\R_DATA_TEMPR0[42] , 
        \Z\R_DATA_TEMPR0[41] , \Z\R_DATA_TEMPR0[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[0][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[0] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[0] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_683 (.A(\Z\R_DATA_TEMPR0[68] ), .B(\Z\R_DATA_TEMPR1[68] ), 
        .C(\Z\R_DATA_TEMPR2[68] ), .D(\Z\R_DATA_TEMPR3[68] ), .Y(
        OR4_683_Y));
    OR4 OR4_209 (.A(\Z\R_DATA_TEMPR16[12] ), .B(\Z\R_DATA_TEMPR17[12] )
        , .C(\Z\R_DATA_TEMPR18[12] ), .D(\Z\R_DATA_TEMPR19[12] ), .Y(
        OR4_209_Y));
    OR4 \OR4_R_DATA[50]  (.A(OR4_131_Y), .B(OR4_300_Y), .C(OR4_632_Y), 
        .D(OR4_349_Y), .Y(R_DATA_c[50]));
    OR4 OR4_516 (.A(\Z\R_DATA_TEMPR8[5] ), .B(\Z\R_DATA_TEMPR9[5] ), 
        .C(\Z\R_DATA_TEMPR10[5] ), .D(\Z\R_DATA_TEMPR11[5] ), .Y(
        OR4_516_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%15%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C1 (
        .A_DOUT({\Z\R_DATA_TEMPR15[79] , \Z\R_DATA_TEMPR15[78] , 
        \Z\R_DATA_TEMPR15[77] , \Z\R_DATA_TEMPR15[76] , 
        \Z\R_DATA_TEMPR15[75] , \Z\R_DATA_TEMPR15[74] , 
        \Z\R_DATA_TEMPR15[73] , \Z\R_DATA_TEMPR15[72] , 
        \Z\R_DATA_TEMPR15[71] , \Z\R_DATA_TEMPR15[70] , 
        \Z\R_DATA_TEMPR15[69] , \Z\R_DATA_TEMPR15[68] , 
        \Z\R_DATA_TEMPR15[67] , \Z\R_DATA_TEMPR15[66] , 
        \Z\R_DATA_TEMPR15[65] , \Z\R_DATA_TEMPR15[64] , 
        \Z\R_DATA_TEMPR15[63] , \Z\R_DATA_TEMPR15[62] , 
        \Z\R_DATA_TEMPR15[61] , \Z\R_DATA_TEMPR15[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR15[59] , \Z\R_DATA_TEMPR15[58] , 
        \Z\R_DATA_TEMPR15[57] , \Z\R_DATA_TEMPR15[56] , 
        \Z\R_DATA_TEMPR15[55] , \Z\R_DATA_TEMPR15[54] , 
        \Z\R_DATA_TEMPR15[53] , \Z\R_DATA_TEMPR15[52] , 
        \Z\R_DATA_TEMPR15[51] , \Z\R_DATA_TEMPR15[50] , 
        \Z\R_DATA_TEMPR15[49] , \Z\R_DATA_TEMPR15[48] , 
        \Z\R_DATA_TEMPR15[47] , \Z\R_DATA_TEMPR15[46] , 
        \Z\R_DATA_TEMPR15[45] , \Z\R_DATA_TEMPR15[44] , 
        \Z\R_DATA_TEMPR15[43] , \Z\R_DATA_TEMPR15[42] , 
        \Z\R_DATA_TEMPR15[41] , \Z\R_DATA_TEMPR15[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[15][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[3] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[3] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%2%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0 (
        .A_DOUT({\Z\R_DATA_TEMPR2[39] , \Z\R_DATA_TEMPR2[38] , 
        \Z\R_DATA_TEMPR2[37] , \Z\R_DATA_TEMPR2[36] , 
        \Z\R_DATA_TEMPR2[35] , \Z\R_DATA_TEMPR2[34] , 
        \Z\R_DATA_TEMPR2[33] , \Z\R_DATA_TEMPR2[32] , 
        \Z\R_DATA_TEMPR2[31] , \Z\R_DATA_TEMPR2[30] , 
        \Z\R_DATA_TEMPR2[29] , \Z\R_DATA_TEMPR2[28] , 
        \Z\R_DATA_TEMPR2[27] , \Z\R_DATA_TEMPR2[26] , 
        \Z\R_DATA_TEMPR2[25] , \Z\R_DATA_TEMPR2[24] , 
        \Z\R_DATA_TEMPR2[23] , \Z\R_DATA_TEMPR2[22] , 
        \Z\R_DATA_TEMPR2[21] , \Z\R_DATA_TEMPR2[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR2[19] , \Z\R_DATA_TEMPR2[18] , 
        \Z\R_DATA_TEMPR2[17] , \Z\R_DATA_TEMPR2[16] , 
        \Z\R_DATA_TEMPR2[15] , \Z\R_DATA_TEMPR2[14] , 
        \Z\R_DATA_TEMPR2[13] , \Z\R_DATA_TEMPR2[12] , 
        \Z\R_DATA_TEMPR2[11] , \Z\R_DATA_TEMPR2[10] , 
        \Z\R_DATA_TEMPR2[9] , \Z\R_DATA_TEMPR2[8] , 
        \Z\R_DATA_TEMPR2[7] , \Z\R_DATA_TEMPR2[6] , 
        \Z\R_DATA_TEMPR2[5] , \Z\R_DATA_TEMPR2[4] , 
        \Z\R_DATA_TEMPR2[3] , \Z\R_DATA_TEMPR2[2] , 
        \Z\R_DATA_TEMPR2[1] , \Z\R_DATA_TEMPR2[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[2][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[0] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[0] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_279 (.A(OR4_436_Y), .B(OR2_66_Y), .C(
        \Z\R_DATA_TEMPR22[56] ), .D(\Z\R_DATA_TEMPR23[56] ), .Y(
        OR4_279_Y));
    OR4 \OR4_R_DATA[63]  (.A(OR4_658_Y), .B(OR4_469_Y), .C(OR4_435_Y), 
        .D(OR4_420_Y), .Y(R_DATA_c[63]));
    OR4 OR4_436 (.A(\Z\R_DATA_TEMPR16[56] ), .B(\Z\R_DATA_TEMPR17[56] )
        , .C(\Z\R_DATA_TEMPR18[56] ), .D(\Z\R_DATA_TEMPR19[56] ), .Y(
        OR4_436_Y));
    OR4 OR4_89 (.A(\Z\R_DATA_TEMPR16[73] ), .B(\Z\R_DATA_TEMPR17[73] ), 
        .C(\Z\R_DATA_TEMPR18[73] ), .D(\Z\R_DATA_TEMPR19[73] ), .Y(
        OR4_89_Y));
    OR4 OR4_453 (.A(\Z\R_DATA_TEMPR4[3] ), .B(\Z\R_DATA_TEMPR5[3] ), 
        .C(\Z\R_DATA_TEMPR6[3] ), .D(\Z\R_DATA_TEMPR7[3] ), .Y(
        OR4_453_Y));
    OR4 \OR4_R_DATA[56]  (.A(OR4_608_Y), .B(OR4_279_Y), .C(OR4_401_Y), 
        .D(OR4_431_Y), .Y(R_DATA_c[56]));
    OR4 OR4_651 (.A(\Z\R_DATA_TEMPR4[50] ), .B(\Z\R_DATA_TEMPR5[50] ), 
        .C(\Z\R_DATA_TEMPR6[50] ), .D(\Z\R_DATA_TEMPR7[50] ), .Y(
        OR4_651_Y));
    OR4 OR4_198 (.A(\Z\R_DATA_TEMPR16[65] ), .B(\Z\R_DATA_TEMPR17[65] )
        , .C(\Z\R_DATA_TEMPR18[65] ), .D(\Z\R_DATA_TEMPR19[65] ), .Y(
        OR4_198_Y));
    OR4 OR4_258 (.A(OR4_587_Y), .B(OR2_16_Y), .C(
        \Z\R_DATA_TEMPR22[48] ), .D(\Z\R_DATA_TEMPR23[48] ), .Y(
        OR4_258_Y));
    OR4 \OR4_R_DATA[21]  (.A(OR4_669_Y), .B(OR4_635_Y), .C(OR4_647_Y), 
        .D(OR4_416_Y), .Y(R_DATA_c[21]));
    OR2 OR2_49 (.A(\Z\R_DATA_TEMPR20[7] ), .B(\Z\R_DATA_TEMPR21[7] ), 
        .Y(OR2_49_Y));
    OR4 OR4_620 (.A(\Z\R_DATA_TEMPR12[43] ), .B(\Z\R_DATA_TEMPR13[43] )
        , .C(\Z\R_DATA_TEMPR14[43] ), .D(\Z\R_DATA_TEMPR15[43] ), .Y(
        OR4_620_Y));
    OR4 OR4_183 (.A(OR4_305_Y), .B(OR4_8_Y), .C(OR4_159_Y), .D(
        OR4_522_Y), .Y(OR4_183_Y));
    OR4 OR4_332 (.A(\Z\R_DATA_TEMPR28[36] ), .B(\Z\R_DATA_TEMPR29[36] )
        , .C(\Z\R_DATA_TEMPR30[36] ), .D(\Z\R_DATA_TEMPR31[36] ), .Y(
        OR4_332_Y));
    OR4 OR4_247 (.A(OR4_106_Y), .B(OR4_276_Y), .C(OR4_346_Y), .D(
        OR4_152_Y), .Y(OR4_247_Y));
    OR4 OR4_13 (.A(\Z\R_DATA_TEMPR28[48] ), .B(\Z\R_DATA_TEMPR29[48] ), 
        .C(\Z\R_DATA_TEMPR30[48] ), .D(\Z\R_DATA_TEMPR31[48] ), .Y(
        OR4_13_Y));
    OR4 OR4_518 (.A(\Z\R_DATA_TEMPR16[40] ), .B(\Z\R_DATA_TEMPR17[40] )
        , .C(\Z\R_DATA_TEMPR18[40] ), .D(\Z\R_DATA_TEMPR19[40] ), .Y(
        OR4_518_Y));
    OR4 OR4_327 (.A(\Z\R_DATA_TEMPR4[6] ), .B(\Z\R_DATA_TEMPR5[6] ), 
        .C(\Z\R_DATA_TEMPR6[6] ), .D(\Z\R_DATA_TEMPR7[6] ), .Y(
        OR4_327_Y));
    OR4 OR4_147 (.A(\Z\R_DATA_TEMPR0[62] ), .B(\Z\R_DATA_TEMPR1[62] ), 
        .C(\Z\R_DATA_TEMPR2[62] ), .D(\Z\R_DATA_TEMPR3[62] ), .Y(
        OR4_147_Y));
    OR4 OR4_120 (.A(\Z\R_DATA_TEMPR28[41] ), .B(\Z\R_DATA_TEMPR29[41] )
        , .C(\Z\R_DATA_TEMPR30[41] ), .D(\Z\R_DATA_TEMPR31[41] ), .Y(
        OR4_120_Y));
    OR4 OR4_51 (.A(\Z\R_DATA_TEMPR8[52] ), .B(\Z\R_DATA_TEMPR9[52] ), 
        .C(\Z\R_DATA_TEMPR10[52] ), .D(\Z\R_DATA_TEMPR11[52] ), .Y(
        OR4_51_Y));
    INV \INVBLKY1[0]  (.A(R_ADDR_c[10]), .Y(\Z\BLKY1[0] ));
    OR2 OR2_2 (.A(\Z\R_DATA_TEMPR20[52] ), .B(\Z\R_DATA_TEMPR21[52] ), 
        .Y(OR2_2_Y));
    OR4 \OR4_R_DATA[20]  (.A(OR4_534_Y), .B(OR4_698_Y), .C(OR4_301_Y), 
        .D(OR4_26_Y), .Y(R_DATA_c[20]));
    CFG2 #( .INIT(4'h8) )  CFG2_5 (.A(R_ADDR_c[12]), .B(R_ADDR_c[11]), 
        .Y(CFG2_5_Y));
    OR2 OR2_69 (.A(\Z\R_DATA_TEMPR20[0] ), .B(\Z\R_DATA_TEMPR21[0] ), 
        .Y(OR2_69_Y));
    OR4 OR4_707 (.A(\Z\R_DATA_TEMPR28[45] ), .B(\Z\R_DATA_TEMPR29[45] )
        , .C(\Z\R_DATA_TEMPR30[45] ), .D(\Z\R_DATA_TEMPR31[45] ), .Y(
        OR4_707_Y));
    OR4 OR4_704 (.A(\Z\R_DATA_TEMPR4[29] ), .B(\Z\R_DATA_TEMPR5[29] ), 
        .C(\Z\R_DATA_TEMPR6[29] ), .D(\Z\R_DATA_TEMPR7[29] ), .Y(
        OR4_704_Y));
    OR4 OR4_20 (.A(\Z\R_DATA_TEMPR8[24] ), .B(\Z\R_DATA_TEMPR9[24] ), 
        .C(\Z\R_DATA_TEMPR10[24] ), .D(\Z\R_DATA_TEMPR11[24] ), .Y(
        OR4_20_Y));
    OR2 OR2_39 (.A(\Z\R_DATA_TEMPR20[31] ), .B(\Z\R_DATA_TEMPR21[31] ), 
        .Y(OR2_39_Y));
    OR4 \OR4_R_DATA[26]  (.A(OR4_280_Y), .B(OR4_673_Y), .C(OR4_68_Y), 
        .D(OR4_101_Y), .Y(R_DATA_c[26]));
    OR4 OR4_416 (.A(\Z\R_DATA_TEMPR28[21] ), .B(\Z\R_DATA_TEMPR29[21] )
        , .C(\Z\R_DATA_TEMPR30[21] ), .D(\Z\R_DATA_TEMPR31[21] ), .Y(
        OR4_416_Y));
    OR4 OR4_244 (.A(\Z\R_DATA_TEMPR12[18] ), .B(\Z\R_DATA_TEMPR13[18] )
        , .C(\Z\R_DATA_TEMPR14[18] ), .D(\Z\R_DATA_TEMPR15[18] ), .Y(
        OR4_244_Y));
    OR4 OR4_27 (.A(\Z\R_DATA_TEMPR24[6] ), .B(\Z\R_DATA_TEMPR25[6] ), 
        .C(\Z\R_DATA_TEMPR26[6] ), .D(\Z\R_DATA_TEMPR27[6] ), .Y(
        OR4_27_Y));
    OR2 OR2_58 (.A(\Z\R_DATA_TEMPR20[37] ), .B(\Z\R_DATA_TEMPR21[37] ), 
        .Y(OR2_58_Y));
    OR4 OR4_82 (.A(\Z\R_DATA_TEMPR12[20] ), .B(\Z\R_DATA_TEMPR13[20] ), 
        .C(\Z\R_DATA_TEMPR14[20] ), .D(\Z\R_DATA_TEMPR15[20] ), .Y(
        OR4_82_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%15%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0 (
        .A_DOUT({\Z\R_DATA_TEMPR15[39] , \Z\R_DATA_TEMPR15[38] , 
        \Z\R_DATA_TEMPR15[37] , \Z\R_DATA_TEMPR15[36] , 
        \Z\R_DATA_TEMPR15[35] , \Z\R_DATA_TEMPR15[34] , 
        \Z\R_DATA_TEMPR15[33] , \Z\R_DATA_TEMPR15[32] , 
        \Z\R_DATA_TEMPR15[31] , \Z\R_DATA_TEMPR15[30] , 
        \Z\R_DATA_TEMPR15[29] , \Z\R_DATA_TEMPR15[28] , 
        \Z\R_DATA_TEMPR15[27] , \Z\R_DATA_TEMPR15[26] , 
        \Z\R_DATA_TEMPR15[25] , \Z\R_DATA_TEMPR15[24] , 
        \Z\R_DATA_TEMPR15[23] , \Z\R_DATA_TEMPR15[22] , 
        \Z\R_DATA_TEMPR15[21] , \Z\R_DATA_TEMPR15[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR15[19] , \Z\R_DATA_TEMPR15[18] , 
        \Z\R_DATA_TEMPR15[17] , \Z\R_DATA_TEMPR15[16] , 
        \Z\R_DATA_TEMPR15[15] , \Z\R_DATA_TEMPR15[14] , 
        \Z\R_DATA_TEMPR15[13] , \Z\R_DATA_TEMPR15[12] , 
        \Z\R_DATA_TEMPR15[11] , \Z\R_DATA_TEMPR15[10] , 
        \Z\R_DATA_TEMPR15[9] , \Z\R_DATA_TEMPR15[8] , 
        \Z\R_DATA_TEMPR15[7] , \Z\R_DATA_TEMPR15[6] , 
        \Z\R_DATA_TEMPR15[5] , \Z\R_DATA_TEMPR15[4] , 
        \Z\R_DATA_TEMPR15[3] , \Z\R_DATA_TEMPR15[2] , 
        \Z\R_DATA_TEMPR15[1] , \Z\R_DATA_TEMPR15[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[15][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[3] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[3] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_230 (.A(OR4_464_Y), .B(OR4_590_Y), .C(OR4_586_Y), .D(
        OR4_710_Y), .Y(OR4_230_Y));
    OR4 OR4_128 (.A(\Z\R_DATA_TEMPR16[22] ), .B(\Z\R_DATA_TEMPR17[22] )
        , .C(\Z\R_DATA_TEMPR18[22] ), .D(\Z\R_DATA_TEMPR19[22] ), .Y(
        OR4_128_Y));
    OR4 OR4_537 (.A(\Z\R_DATA_TEMPR4[68] ), .B(\Z\R_DATA_TEMPR5[68] ), 
        .C(\Z\R_DATA_TEMPR6[68] ), .D(\Z\R_DATA_TEMPR7[68] ), .Y(
        OR4_537_Y));
    OR2 OR2_42 (.A(\Z\R_DATA_TEMPR20[8] ), .B(\Z\R_DATA_TEMPR21[8] ), 
        .Y(OR2_42_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%17%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0 (
        .A_DOUT({\Z\R_DATA_TEMPR17[39] , \Z\R_DATA_TEMPR17[38] , 
        \Z\R_DATA_TEMPR17[37] , \Z\R_DATA_TEMPR17[36] , 
        \Z\R_DATA_TEMPR17[35] , \Z\R_DATA_TEMPR17[34] , 
        \Z\R_DATA_TEMPR17[33] , \Z\R_DATA_TEMPR17[32] , 
        \Z\R_DATA_TEMPR17[31] , \Z\R_DATA_TEMPR17[30] , 
        \Z\R_DATA_TEMPR17[29] , \Z\R_DATA_TEMPR17[28] , 
        \Z\R_DATA_TEMPR17[27] , \Z\R_DATA_TEMPR17[26] , 
        \Z\R_DATA_TEMPR17[25] , \Z\R_DATA_TEMPR17[24] , 
        \Z\R_DATA_TEMPR17[23] , \Z\R_DATA_TEMPR17[22] , 
        \Z\R_DATA_TEMPR17[21] , \Z\R_DATA_TEMPR17[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR17[19] , \Z\R_DATA_TEMPR17[18] , 
        \Z\R_DATA_TEMPR17[17] , \Z\R_DATA_TEMPR17[16] , 
        \Z\R_DATA_TEMPR17[15] , \Z\R_DATA_TEMPR17[14] , 
        \Z\R_DATA_TEMPR17[13] , \Z\R_DATA_TEMPR17[12] , 
        \Z\R_DATA_TEMPR17[11] , \Z\R_DATA_TEMPR17[10] , 
        \Z\R_DATA_TEMPR17[9] , \Z\R_DATA_TEMPR17[8] , 
        \Z\R_DATA_TEMPR17[7] , \Z\R_DATA_TEMPR17[6] , 
        \Z\R_DATA_TEMPR17[5] , \Z\R_DATA_TEMPR17[4] , 
        \Z\R_DATA_TEMPR17[3] , \Z\R_DATA_TEMPR17[2] , 
        \Z\R_DATA_TEMPR17[1] , \Z\R_DATA_TEMPR17[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[17][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[4] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[4] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_182 (.A(\Z\R_DATA_TEMPR16[16] ), .B(\Z\R_DATA_TEMPR17[16] )
        , .C(\Z\R_DATA_TEMPR18[16] ), .D(\Z\R_DATA_TEMPR19[16] ), .Y(
        OR4_182_Y));
    OR4 OR4_465 (.A(\Z\R_DATA_TEMPR8[58] ), .B(\Z\R_DATA_TEMPR9[58] ), 
        .C(\Z\R_DATA_TEMPR10[58] ), .D(\Z\R_DATA_TEMPR11[58] ), .Y(
        OR4_465_Y));
    OR4 OR4_312 (.A(\Z\R_DATA_TEMPR28[4] ), .B(\Z\R_DATA_TEMPR29[4] ), 
        .C(\Z\R_DATA_TEMPR30[4] ), .D(\Z\R_DATA_TEMPR31[4] ), .Y(
        OR4_312_Y));
    OR4 OR4_64 (.A(\Z\R_DATA_TEMPR8[53] ), .B(\Z\R_DATA_TEMPR9[53] ), 
        .C(\Z\R_DATA_TEMPR10[53] ), .D(\Z\R_DATA_TEMPR11[53] ), .Y(
        OR4_64_Y));
    OR4 OR4_551 (.A(\Z\R_DATA_TEMPR28[2] ), .B(\Z\R_DATA_TEMPR29[2] ), 
        .C(\Z\R_DATA_TEMPR30[2] ), .D(\Z\R_DATA_TEMPR31[2] ), .Y(
        OR4_551_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%23%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C1 (
        .A_DOUT({\Z\R_DATA_TEMPR23[79] , \Z\R_DATA_TEMPR23[78] , 
        \Z\R_DATA_TEMPR23[77] , \Z\R_DATA_TEMPR23[76] , 
        \Z\R_DATA_TEMPR23[75] , \Z\R_DATA_TEMPR23[74] , 
        \Z\R_DATA_TEMPR23[73] , \Z\R_DATA_TEMPR23[72] , 
        \Z\R_DATA_TEMPR23[71] , \Z\R_DATA_TEMPR23[70] , 
        \Z\R_DATA_TEMPR23[69] , \Z\R_DATA_TEMPR23[68] , 
        \Z\R_DATA_TEMPR23[67] , \Z\R_DATA_TEMPR23[66] , 
        \Z\R_DATA_TEMPR23[65] , \Z\R_DATA_TEMPR23[64] , 
        \Z\R_DATA_TEMPR23[63] , \Z\R_DATA_TEMPR23[62] , 
        \Z\R_DATA_TEMPR23[61] , \Z\R_DATA_TEMPR23[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR23[59] , \Z\R_DATA_TEMPR23[58] , 
        \Z\R_DATA_TEMPR23[57] , \Z\R_DATA_TEMPR23[56] , 
        \Z\R_DATA_TEMPR23[55] , \Z\R_DATA_TEMPR23[54] , 
        \Z\R_DATA_TEMPR23[53] , \Z\R_DATA_TEMPR23[52] , 
        \Z\R_DATA_TEMPR23[51] , \Z\R_DATA_TEMPR23[50] , 
        \Z\R_DATA_TEMPR23[49] , \Z\R_DATA_TEMPR23[48] , 
        \Z\R_DATA_TEMPR23[47] , \Z\R_DATA_TEMPR23[46] , 
        \Z\R_DATA_TEMPR23[45] , \Z\R_DATA_TEMPR23[44] , 
        \Z\R_DATA_TEMPR23[43] , \Z\R_DATA_TEMPR23[42] , 
        \Z\R_DATA_TEMPR23[41] , \Z\R_DATA_TEMPR23[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[23][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[5] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[5] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_11 (.A(\Z\R_DATA_TEMPR4[1] ), .B(\Z\R_DATA_TEMPR5[1] ), .C(
        \Z\R_DATA_TEMPR6[1] ), .D(\Z\R_DATA_TEMPR7[1] ), .Y(OR4_11_Y));
    OR4 OR4_639 (.A(\Z\R_DATA_TEMPR4[9] ), .B(\Z\R_DATA_TEMPR5[9] ), 
        .C(\Z\R_DATA_TEMPR6[9] ), .D(\Z\R_DATA_TEMPR7[9] ), .Y(
        OR4_639_Y));
    OR4 OR4_345 (.A(\Z\R_DATA_TEMPR16[31] ), .B(\Z\R_DATA_TEMPR17[31] )
        , .C(\Z\R_DATA_TEMPR18[31] ), .D(\Z\R_DATA_TEMPR19[31] ), .Y(
        OR4_345_Y));
    OR4 OR4_236 (.A(\Z\R_DATA_TEMPR24[13] ), .B(\Z\R_DATA_TEMPR25[13] )
        , .C(\Z\R_DATA_TEMPR26[13] ), .D(\Z\R_DATA_TEMPR27[13] ), .Y(
        OR4_236_Y));
    OR2 OR2_7 (.A(\Z\R_DATA_TEMPR20[69] ), .B(\Z\R_DATA_TEMPR21[69] ), 
        .Y(OR2_7_Y));
    OR4 OR4_73 (.A(\Z\R_DATA_TEMPR12[36] ), .B(\Z\R_DATA_TEMPR13[36] ), 
        .C(\Z\R_DATA_TEMPR14[36] ), .D(\Z\R_DATA_TEMPR15[36] ), .Y(
        OR4_73_Y));
    OR4 OR4_195 (.A(\Z\R_DATA_TEMPR0[77] ), .B(\Z\R_DATA_TEMPR1[77] ), 
        .C(\Z\R_DATA_TEMPR2[77] ), .D(\Z\R_DATA_TEMPR3[77] ), .Y(
        OR4_195_Y));
    OR2 OR2_62 (.A(\Z\R_DATA_TEMPR20[4] ), .B(\Z\R_DATA_TEMPR21[4] ), 
        .Y(OR2_62_Y));
    OR4 OR4_252 (.A(OR4_555_Y), .B(OR2_65_Y), .C(
        \Z\R_DATA_TEMPR22[39] ), .D(\Z\R_DATA_TEMPR23[39] ), .Y(
        OR4_252_Y));
    OR4 OR4_289 (.A(\Z\R_DATA_TEMPR4[78] ), .B(\Z\R_DATA_TEMPR5[78] ), 
        .C(\Z\R_DATA_TEMPR6[78] ), .D(\Z\R_DATA_TEMPR7[78] ), .Y(
        OR4_289_Y));
    OR4 OR4_497 (.A(OR4_61_Y), .B(OR4_304_Y), .C(OR4_619_Y), .D(
        OR4_203_Y), .Y(OR4_497_Y));
    OR2 OR2_32 (.A(\Z\R_DATA_TEMPR20[11] ), .B(\Z\R_DATA_TEMPR21[11] ), 
        .Y(OR2_32_Y));
    OR4 OR4_634 (.A(\Z\R_DATA_TEMPR28[58] ), .B(\Z\R_DATA_TEMPR29[58] )
        , .C(\Z\R_DATA_TEMPR30[58] ), .D(\Z\R_DATA_TEMPR31[58] ), .Y(
        OR4_634_Y));
    OR2 OR2_1 (.A(\Z\R_DATA_TEMPR20[78] ), .B(\Z\R_DATA_TEMPR21[78] ), 
        .Y(OR2_1_Y));
    OR4 OR4_464 (.A(\Z\R_DATA_TEMPR0[61] ), .B(\Z\R_DATA_TEMPR1[61] ), 
        .C(\Z\R_DATA_TEMPR2[61] ), .D(\Z\R_DATA_TEMPR3[61] ), .Y(
        OR4_464_Y));
    OR4 \OR4_R_DATA[57]  (.A(OR4_421_Y), .B(OR4_43_Y), .C(OR4_241_Y), 
        .D(OR4_294_Y), .Y(R_DATA_c[57]));
    OR4 OR4_210 (.A(\Z\R_DATA_TEMPR24[61] ), .B(\Z\R_DATA_TEMPR25[61] )
        , .C(\Z\R_DATA_TEMPR26[61] ), .D(\Z\R_DATA_TEMPR27[61] ), .Y(
        OR4_210_Y));
    OR4 OR4_517 (.A(\Z\R_DATA_TEMPR0[51] ), .B(\Z\R_DATA_TEMPR1[51] ), 
        .C(\Z\R_DATA_TEMPR2[51] ), .D(\Z\R_DATA_TEMPR3[51] ), .Y(
        OR4_517_Y));
    OR4 OR4_350 (.A(\Z\R_DATA_TEMPR24[66] ), .B(\Z\R_DATA_TEMPR25[66] )
        , .C(\Z\R_DATA_TEMPR26[66] ), .D(\Z\R_DATA_TEMPR27[66] ), .Y(
        OR4_350_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%31%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C1 (
        .A_DOUT({\Z\R_DATA_TEMPR31[79] , \Z\R_DATA_TEMPR31[78] , 
        \Z\R_DATA_TEMPR31[77] , \Z\R_DATA_TEMPR31[76] , 
        \Z\R_DATA_TEMPR31[75] , \Z\R_DATA_TEMPR31[74] , 
        \Z\R_DATA_TEMPR31[73] , \Z\R_DATA_TEMPR31[72] , 
        \Z\R_DATA_TEMPR31[71] , \Z\R_DATA_TEMPR31[70] , 
        \Z\R_DATA_TEMPR31[69] , \Z\R_DATA_TEMPR31[68] , 
        \Z\R_DATA_TEMPR31[67] , \Z\R_DATA_TEMPR31[66] , 
        \Z\R_DATA_TEMPR31[65] , \Z\R_DATA_TEMPR31[64] , 
        \Z\R_DATA_TEMPR31[63] , \Z\R_DATA_TEMPR31[62] , 
        \Z\R_DATA_TEMPR31[61] , \Z\R_DATA_TEMPR31[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR31[59] , \Z\R_DATA_TEMPR31[58] , 
        \Z\R_DATA_TEMPR31[57] , \Z\R_DATA_TEMPR31[56] , 
        \Z\R_DATA_TEMPR31[55] , \Z\R_DATA_TEMPR31[54] , 
        \Z\R_DATA_TEMPR31[53] , \Z\R_DATA_TEMPR31[52] , 
        \Z\R_DATA_TEMPR31[51] , \Z\R_DATA_TEMPR31[50] , 
        \Z\R_DATA_TEMPR31[49] , \Z\R_DATA_TEMPR31[48] , 
        \Z\R_DATA_TEMPR31[47] , \Z\R_DATA_TEMPR31[46] , 
        \Z\R_DATA_TEMPR31[45] , \Z\R_DATA_TEMPR31[44] , 
        \Z\R_DATA_TEMPR31[43] , \Z\R_DATA_TEMPR31[42] , 
        \Z\R_DATA_TEMPR31[41] , \Z\R_DATA_TEMPR31[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[31][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[7] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[7] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%24%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0 (
        .A_DOUT({\Z\R_DATA_TEMPR24[39] , \Z\R_DATA_TEMPR24[38] , 
        \Z\R_DATA_TEMPR24[37] , \Z\R_DATA_TEMPR24[36] , 
        \Z\R_DATA_TEMPR24[35] , \Z\R_DATA_TEMPR24[34] , 
        \Z\R_DATA_TEMPR24[33] , \Z\R_DATA_TEMPR24[32] , 
        \Z\R_DATA_TEMPR24[31] , \Z\R_DATA_TEMPR24[30] , 
        \Z\R_DATA_TEMPR24[29] , \Z\R_DATA_TEMPR24[28] , 
        \Z\R_DATA_TEMPR24[27] , \Z\R_DATA_TEMPR24[26] , 
        \Z\R_DATA_TEMPR24[25] , \Z\R_DATA_TEMPR24[24] , 
        \Z\R_DATA_TEMPR24[23] , \Z\R_DATA_TEMPR24[22] , 
        \Z\R_DATA_TEMPR24[21] , \Z\R_DATA_TEMPR24[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR24[19] , \Z\R_DATA_TEMPR24[18] , 
        \Z\R_DATA_TEMPR24[17] , \Z\R_DATA_TEMPR24[16] , 
        \Z\R_DATA_TEMPR24[15] , \Z\R_DATA_TEMPR24[14] , 
        \Z\R_DATA_TEMPR24[13] , \Z\R_DATA_TEMPR24[12] , 
        \Z\R_DATA_TEMPR24[11] , \Z\R_DATA_TEMPR24[10] , 
        \Z\R_DATA_TEMPR24[9] , \Z\R_DATA_TEMPR24[8] , 
        \Z\R_DATA_TEMPR24[7] , \Z\R_DATA_TEMPR24[6] , 
        \Z\R_DATA_TEMPR24[5] , \Z\R_DATA_TEMPR24[4] , 
        \Z\R_DATA_TEMPR24[3] , \Z\R_DATA_TEMPR24[2] , 
        \Z\R_DATA_TEMPR24[1] , \Z\R_DATA_TEMPR24[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[24][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[6] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[6] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_366 (.A(\Z\R_DATA_TEMPR28[33] ), .B(\Z\R_DATA_TEMPR29[33] )
        , .C(\Z\R_DATA_TEMPR30[33] ), .D(\Z\R_DATA_TEMPR31[33] ), .Y(
        OR4_366_Y));
    OR4 OR4_295 (.A(\Z\R_DATA_TEMPR8[64] ), .B(\Z\R_DATA_TEMPR9[64] ), 
        .C(\Z\R_DATA_TEMPR10[64] ), .D(\Z\R_DATA_TEMPR11[64] ), .Y(
        OR4_295_Y));
    OR4 \OR4_R_DATA[72]  (.A(OR4_495_Y), .B(OR4_476_Y), .C(OR4_372_Y), 
        .D(OR4_45_Y), .Y(R_DATA_c[72]));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%19%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C1 (
        .A_DOUT({\Z\R_DATA_TEMPR19[79] , \Z\R_DATA_TEMPR19[78] , 
        \Z\R_DATA_TEMPR19[77] , \Z\R_DATA_TEMPR19[76] , 
        \Z\R_DATA_TEMPR19[75] , \Z\R_DATA_TEMPR19[74] , 
        \Z\R_DATA_TEMPR19[73] , \Z\R_DATA_TEMPR19[72] , 
        \Z\R_DATA_TEMPR19[71] , \Z\R_DATA_TEMPR19[70] , 
        \Z\R_DATA_TEMPR19[69] , \Z\R_DATA_TEMPR19[68] , 
        \Z\R_DATA_TEMPR19[67] , \Z\R_DATA_TEMPR19[66] , 
        \Z\R_DATA_TEMPR19[65] , \Z\R_DATA_TEMPR19[64] , 
        \Z\R_DATA_TEMPR19[63] , \Z\R_DATA_TEMPR19[62] , 
        \Z\R_DATA_TEMPR19[61] , \Z\R_DATA_TEMPR19[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR19[59] , \Z\R_DATA_TEMPR19[58] , 
        \Z\R_DATA_TEMPR19[57] , \Z\R_DATA_TEMPR19[56] , 
        \Z\R_DATA_TEMPR19[55] , \Z\R_DATA_TEMPR19[54] , 
        \Z\R_DATA_TEMPR19[53] , \Z\R_DATA_TEMPR19[52] , 
        \Z\R_DATA_TEMPR19[51] , \Z\R_DATA_TEMPR19[50] , 
        \Z\R_DATA_TEMPR19[49] , \Z\R_DATA_TEMPR19[48] , 
        \Z\R_DATA_TEMPR19[47] , \Z\R_DATA_TEMPR19[46] , 
        \Z\R_DATA_TEMPR19[45] , \Z\R_DATA_TEMPR19[44] , 
        \Z\R_DATA_TEMPR19[43] , \Z\R_DATA_TEMPR19[42] , 
        \Z\R_DATA_TEMPR19[41] , \Z\R_DATA_TEMPR19[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[19][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[4] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[4] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_645 (.A(\Z\R_DATA_TEMPR12[16] ), .B(\Z\R_DATA_TEMPR13[16] )
        , .C(\Z\R_DATA_TEMPR14[16] ), .D(\Z\R_DATA_TEMPR15[16] ), .Y(
        OR4_645_Y));
    OR4 OR4_619 (.A(\Z\R_DATA_TEMPR8[59] ), .B(\Z\R_DATA_TEMPR9[59] ), 
        .C(\Z\R_DATA_TEMPR10[59] ), .D(\Z\R_DATA_TEMPR11[59] ), .Y(
        OR4_619_Y));
    OR4 OR4_35 (.A(\Z\R_DATA_TEMPR4[40] ), .B(\Z\R_DATA_TEMPR5[40] ), 
        .C(\Z\R_DATA_TEMPR6[40] ), .D(\Z\R_DATA_TEMPR7[40] ), .Y(
        OR4_35_Y));
    OR4 OR4_405 (.A(\Z\R_DATA_TEMPR0[28] ), .B(\Z\R_DATA_TEMPR1[28] ), 
        .C(\Z\R_DATA_TEMPR2[28] ), .D(\Z\R_DATA_TEMPR3[28] ), .Y(
        OR4_405_Y));
    OR4 OR4_216 (.A(\Z\R_DATA_TEMPR0[52] ), .B(\Z\R_DATA_TEMPR1[52] ), 
        .C(\Z\R_DATA_TEMPR2[52] ), .D(\Z\R_DATA_TEMPR3[52] ), .Y(
        OR4_216_Y));
    OR4 OR4_71 (.A(\Z\R_DATA_TEMPR8[14] ), .B(\Z\R_DATA_TEMPR9[14] ), 
        .C(\Z\R_DATA_TEMPR10[14] ), .D(\Z\R_DATA_TEMPR11[14] ), .Y(
        OR4_71_Y));
    OR4 OR4_475 (.A(\Z\R_DATA_TEMPR0[20] ), .B(\Z\R_DATA_TEMPR1[20] ), 
        .C(\Z\R_DATA_TEMPR2[20] ), .D(\Z\R_DATA_TEMPR3[20] ), .Y(
        OR4_475_Y));
    OR4 OR4_125 (.A(OR4_638_Y), .B(OR4_488_Y), .C(OR4_365_Y), .D(
        OR4_396_Y), .Y(OR4_125_Y));
    OR4 OR4_493 (.A(\Z\R_DATA_TEMPR24[53] ), .B(\Z\R_DATA_TEMPR25[53] )
        , .C(\Z\R_DATA_TEMPR26[53] ), .D(\Z\R_DATA_TEMPR27[53] ), .Y(
        OR4_493_Y));
    OR4 OR4_691 (.A(OR4_187_Y), .B(OR2_32_Y), .C(
        \Z\R_DATA_TEMPR22[11] ), .D(\Z\R_DATA_TEMPR23[11] ), .Y(
        OR4_691_Y));
    OR4 OR4_614 (.A(\Z\R_DATA_TEMPR4[17] ), .B(\Z\R_DATA_TEMPR5[17] ), 
        .C(\Z\R_DATA_TEMPR6[17] ), .D(\Z\R_DATA_TEMPR7[17] ), .Y(
        OR4_614_Y));
    OR4 OR4_427 (.A(\Z\R_DATA_TEMPR16[1] ), .B(\Z\R_DATA_TEMPR17[1] ), 
        .C(\Z\R_DATA_TEMPR18[1] ), .D(\Z\R_DATA_TEMPR19[1] ), .Y(
        OR4_427_Y));
    OR4 OR4_298 (.A(\Z\R_DATA_TEMPR28[75] ), .B(\Z\R_DATA_TEMPR29[75] )
        , .C(\Z\R_DATA_TEMPR30[75] ), .D(\Z\R_DATA_TEMPR31[75] ), .Y(
        OR4_298_Y));
    OR4 \OR4_R_DATA[27]  (.A(OR4_87_Y), .B(OR4_433_Y), .C(OR4_624_Y), 
        .D(OR4_692_Y), .Y(R_DATA_c[27]));
    OR4 OR4_28 (.A(\Z\R_DATA_TEMPR24[65] ), .B(\Z\R_DATA_TEMPR25[65] ), 
        .C(\Z\R_DATA_TEMPR26[65] ), .D(\Z\R_DATA_TEMPR27[65] ), .Y(
        OR4_28_Y));
    OR4 OR4_640 (.A(\Z\R_DATA_TEMPR8[51] ), .B(\Z\R_DATA_TEMPR9[51] ), 
        .C(\Z\R_DATA_TEMPR10[51] ), .D(\Z\R_DATA_TEMPR11[51] ), .Y(
        OR4_640_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%8%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0 (
        .A_DOUT({\Z\R_DATA_TEMPR8[39] , \Z\R_DATA_TEMPR8[38] , 
        \Z\R_DATA_TEMPR8[37] , \Z\R_DATA_TEMPR8[36] , 
        \Z\R_DATA_TEMPR8[35] , \Z\R_DATA_TEMPR8[34] , 
        \Z\R_DATA_TEMPR8[33] , \Z\R_DATA_TEMPR8[32] , 
        \Z\R_DATA_TEMPR8[31] , \Z\R_DATA_TEMPR8[30] , 
        \Z\R_DATA_TEMPR8[29] , \Z\R_DATA_TEMPR8[28] , 
        \Z\R_DATA_TEMPR8[27] , \Z\R_DATA_TEMPR8[26] , 
        \Z\R_DATA_TEMPR8[25] , \Z\R_DATA_TEMPR8[24] , 
        \Z\R_DATA_TEMPR8[23] , \Z\R_DATA_TEMPR8[22] , 
        \Z\R_DATA_TEMPR8[21] , \Z\R_DATA_TEMPR8[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR8[19] , \Z\R_DATA_TEMPR8[18] , 
        \Z\R_DATA_TEMPR8[17] , \Z\R_DATA_TEMPR8[16] , 
        \Z\R_DATA_TEMPR8[15] , \Z\R_DATA_TEMPR8[14] , 
        \Z\R_DATA_TEMPR8[13] , \Z\R_DATA_TEMPR8[12] , 
        \Z\R_DATA_TEMPR8[11] , \Z\R_DATA_TEMPR8[10] , 
        \Z\R_DATA_TEMPR8[9] , \Z\R_DATA_TEMPR8[8] , 
        \Z\R_DATA_TEMPR8[7] , \Z\R_DATA_TEMPR8[6] , 
        \Z\R_DATA_TEMPR8[5] , \Z\R_DATA_TEMPR8[4] , 
        \Z\R_DATA_TEMPR8[3] , \Z\R_DATA_TEMPR8[2] , 
        \Z\R_DATA_TEMPR8[1] , \Z\R_DATA_TEMPR8[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[8][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[2] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[2] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[73]  (.A(OR4_412_Y), .B(OR4_235_Y), .C(OR4_213_Y), 
        .D(OR4_180_Y), .Y(R_DATA_c[73]));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKY2[6]  (.A(CFG2_1_Y), .B(
        R_ADDR_c[13]), .C(R_EN_c), .Y(\Z\BLKY2[6] ));
    OR4 OR4_164 (.A(\Z\R_DATA_TEMPR24[23] ), .B(\Z\R_DATA_TEMPR25[23] )
        , .C(\Z\R_DATA_TEMPR26[23] ), .D(\Z\R_DATA_TEMPR27[23] ), .Y(
        OR4_164_Y));
    OR4 OR4_404 (.A(\Z\R_DATA_TEMPR0[65] ), .B(\Z\R_DATA_TEMPR1[65] ), 
        .C(\Z\R_DATA_TEMPR2[65] ), .D(\Z\R_DATA_TEMPR3[65] ), .Y(
        OR4_404_Y));
    OR4 OR4_225 (.A(\Z\R_DATA_TEMPR4[4] ), .B(\Z\R_DATA_TEMPR5[4] ), 
        .C(\Z\R_DATA_TEMPR6[4] ), .D(\Z\R_DATA_TEMPR7[4] ), .Y(
        OR4_225_Y));
    CFG2 #( .INIT(4'h4) )  CFG2_2 (.A(W_ADDR_c[12]), .B(W_ADDR_c[11]), 
        .Y(CFG2_2_Y));
    OR4 OR4_555 (.A(\Z\R_DATA_TEMPR16[39] ), .B(\Z\R_DATA_TEMPR17[39] )
        , .C(\Z\R_DATA_TEMPR18[39] ), .D(\Z\R_DATA_TEMPR19[39] ), .Y(
        OR4_555_Y));
    OR4 OR4_347 (.A(\Z\R_DATA_TEMPR8[19] ), .B(\Z\R_DATA_TEMPR9[19] ), 
        .C(\Z\R_DATA_TEMPR10[19] ), .D(\Z\R_DATA_TEMPR11[19] ), .Y(
        OR4_347_Y));
    OR4 OR4_140 (.A(\Z\R_DATA_TEMPR16[6] ), .B(\Z\R_DATA_TEMPR17[6] ), 
        .C(\Z\R_DATA_TEMPR18[6] ), .D(\Z\R_DATA_TEMPR19[6] ), .Y(
        OR4_140_Y));
    OR4 OR4_474 (.A(\Z\R_DATA_TEMPR0[2] ), .B(\Z\R_DATA_TEMPR1[2] ), 
        .C(\Z\R_DATA_TEMPR2[2] ), .D(\Z\R_DATA_TEMPR3[2] ), .Y(
        OR4_474_Y));
    OR4 OR4_306 (.A(\Z\R_DATA_TEMPR16[30] ), .B(\Z\R_DATA_TEMPR17[30] )
        , .C(\Z\R_DATA_TEMPR18[30] ), .D(\Z\R_DATA_TEMPR19[30] ), .Y(
        OR4_306_Y));
    OR4 OR4_653 (.A(\Z\R_DATA_TEMPR12[31] ), .B(\Z\R_DATA_TEMPR13[31] )
        , .C(\Z\R_DATA_TEMPR14[31] ), .D(\Z\R_DATA_TEMPR15[31] ), .Y(
        OR4_653_Y));
    CFG2 #( .INIT(4'h1) )  CFG2_3 (.A(R_ADDR_c[12]), .B(R_ADDR_c[11]), 
        .Y(CFG2_3_Y));
    OR4 OR4_376 (.A(\Z\R_DATA_TEMPR4[44] ), .B(\Z\R_DATA_TEMPR5[44] ), 
        .C(\Z\R_DATA_TEMPR6[44] ), .D(\Z\R_DATA_TEMPR7[44] ), .Y(
        OR4_376_Y));
    OR4 OR4_423 (.A(\Z\R_DATA_TEMPR12[21] ), .B(\Z\R_DATA_TEMPR13[21] )
        , .C(\Z\R_DATA_TEMPR14[21] ), .D(\Z\R_DATA_TEMPR15[21] ), .Y(
        OR4_423_Y));
    OR4 OR4_84 (.A(OR4_281_Y), .B(OR2_15_Y), .C(\Z\R_DATA_TEMPR22[44] )
        , .D(\Z\R_DATA_TEMPR23[44] ), .Y(OR4_84_Y));
    OR4 OR4_621 (.A(\Z\R_DATA_TEMPR28[19] ), .B(\Z\R_DATA_TEMPR29[19] )
        , .C(\Z\R_DATA_TEMPR30[19] ), .D(\Z\R_DATA_TEMPR31[19] ), .Y(
        OR4_621_Y));
    OR4 OR4_148 (.A(\Z\R_DATA_TEMPR16[28] ), .B(\Z\R_DATA_TEMPR17[28] )
        , .C(\Z\R_DATA_TEMPR18[28] ), .D(\Z\R_DATA_TEMPR19[28] ), .Y(
        OR4_148_Y));
    OR4 OR4_228 (.A(\Z\R_DATA_TEMPR12[5] ), .B(\Z\R_DATA_TEMPR13[5] ), 
        .C(\Z\R_DATA_TEMPR14[5] ), .D(\Z\R_DATA_TEMPR15[5] ), .Y(
        OR4_228_Y));
    OR2 OR2_44 (.A(\Z\R_DATA_TEMPR20[25] ), .B(\Z\R_DATA_TEMPR21[25] ), 
        .Y(OR2_44_Y));
    OR4 OR4_566 (.A(\Z\R_DATA_TEMPR8[69] ), .B(\Z\R_DATA_TEMPR9[69] ), 
        .C(\Z\R_DATA_TEMPR10[69] ), .D(\Z\R_DATA_TEMPR11[69] ), .Y(
        OR4_566_Y));
    OR4 OR4_591 (.A(\Z\R_DATA_TEMPR0[47] ), .B(\Z\R_DATA_TEMPR1[47] ), 
        .C(\Z\R_DATA_TEMPR2[47] ), .D(\Z\R_DATA_TEMPR3[47] ), .Y(
        OR4_591_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%22%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0 (
        .A_DOUT({\Z\R_DATA_TEMPR22[39] , \Z\R_DATA_TEMPR22[38] , 
        \Z\R_DATA_TEMPR22[37] , \Z\R_DATA_TEMPR22[36] , 
        \Z\R_DATA_TEMPR22[35] , \Z\R_DATA_TEMPR22[34] , 
        \Z\R_DATA_TEMPR22[33] , \Z\R_DATA_TEMPR22[32] , 
        \Z\R_DATA_TEMPR22[31] , \Z\R_DATA_TEMPR22[30] , 
        \Z\R_DATA_TEMPR22[29] , \Z\R_DATA_TEMPR22[28] , 
        \Z\R_DATA_TEMPR22[27] , \Z\R_DATA_TEMPR22[26] , 
        \Z\R_DATA_TEMPR22[25] , \Z\R_DATA_TEMPR22[24] , 
        \Z\R_DATA_TEMPR22[23] , \Z\R_DATA_TEMPR22[22] , 
        \Z\R_DATA_TEMPR22[21] , \Z\R_DATA_TEMPR22[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR22[19] , \Z\R_DATA_TEMPR22[18] , 
        \Z\R_DATA_TEMPR22[17] , \Z\R_DATA_TEMPR22[16] , 
        \Z\R_DATA_TEMPR22[15] , \Z\R_DATA_TEMPR22[14] , 
        \Z\R_DATA_TEMPR22[13] , \Z\R_DATA_TEMPR22[12] , 
        \Z\R_DATA_TEMPR22[11] , \Z\R_DATA_TEMPR22[10] , 
        \Z\R_DATA_TEMPR22[9] , \Z\R_DATA_TEMPR22[8] , 
        \Z\R_DATA_TEMPR22[7] , \Z\R_DATA_TEMPR22[6] , 
        \Z\R_DATA_TEMPR22[5] , \Z\R_DATA_TEMPR22[4] , 
        \Z\R_DATA_TEMPR22[3] , \Z\R_DATA_TEMPR22[2] , 
        \Z\R_DATA_TEMPR22[1] , \Z\R_DATA_TEMPR22[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[22][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[5] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[5] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_153 (.A(OR4_46_Y), .B(OR2_38_Y), .C(\Z\R_DATA_TEMPR22[47] )
        , .D(\Z\R_DATA_TEMPR23[47] ), .Y(OR4_153_Y));
    OR4 OR4_9 (.A(OR4_319_Y), .B(OR2_79_Y), .C(\Z\R_DATA_TEMPR22[29] ), 
        .D(\Z\R_DATA_TEMPR23[29] ), .Y(OR4_9_Y));
    OR4 OR4_231 (.A(\Z\R_DATA_TEMPR4[2] ), .B(\Z\R_DATA_TEMPR5[2] ), 
        .C(\Z\R_DATA_TEMPR6[2] ), .D(\Z\R_DATA_TEMPR7[2] ), .Y(
        OR4_231_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%4%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0 (
        .A_DOUT({\Z\R_DATA_TEMPR4[39] , \Z\R_DATA_TEMPR4[38] , 
        \Z\R_DATA_TEMPR4[37] , \Z\R_DATA_TEMPR4[36] , 
        \Z\R_DATA_TEMPR4[35] , \Z\R_DATA_TEMPR4[34] , 
        \Z\R_DATA_TEMPR4[33] , \Z\R_DATA_TEMPR4[32] , 
        \Z\R_DATA_TEMPR4[31] , \Z\R_DATA_TEMPR4[30] , 
        \Z\R_DATA_TEMPR4[29] , \Z\R_DATA_TEMPR4[28] , 
        \Z\R_DATA_TEMPR4[27] , \Z\R_DATA_TEMPR4[26] , 
        \Z\R_DATA_TEMPR4[25] , \Z\R_DATA_TEMPR4[24] , 
        \Z\R_DATA_TEMPR4[23] , \Z\R_DATA_TEMPR4[22] , 
        \Z\R_DATA_TEMPR4[21] , \Z\R_DATA_TEMPR4[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR4[19] , \Z\R_DATA_TEMPR4[18] , 
        \Z\R_DATA_TEMPR4[17] , \Z\R_DATA_TEMPR4[16] , 
        \Z\R_DATA_TEMPR4[15] , \Z\R_DATA_TEMPR4[14] , 
        \Z\R_DATA_TEMPR4[13] , \Z\R_DATA_TEMPR4[12] , 
        \Z\R_DATA_TEMPR4[11] , \Z\R_DATA_TEMPR4[10] , 
        \Z\R_DATA_TEMPR4[9] , \Z\R_DATA_TEMPR4[8] , 
        \Z\R_DATA_TEMPR4[7] , \Z\R_DATA_TEMPR4[6] , 
        \Z\R_DATA_TEMPR4[5] , \Z\R_DATA_TEMPR4[4] , 
        \Z\R_DATA_TEMPR4[3] , \Z\R_DATA_TEMPR4[2] , 
        \Z\R_DATA_TEMPR4[1] , \Z\R_DATA_TEMPR4[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[4][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[1] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[1] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_104 (.A(\Z\R_DATA_TEMPR16[26] ), .B(\Z\R_DATA_TEMPR17[26] )
        , .C(\Z\R_DATA_TEMPR18[26] ), .D(\Z\R_DATA_TEMPR19[26] ), .Y(
        OR4_104_Y));
    OR4 OR4_292 (.A(\Z\R_DATA_TEMPR28[62] ), .B(\Z\R_DATA_TEMPR29[62] )
        , .C(\Z\R_DATA_TEMPR30[62] ), .D(\Z\R_DATA_TEMPR31[62] ), .Y(
        OR4_292_Y));
    OR2 OR2_64 (.A(\Z\R_DATA_TEMPR20[72] ), .B(\Z\R_DATA_TEMPR21[72] ), 
        .Y(OR2_64_Y));
    OR4 OR4_174 (.A(\Z\R_DATA_TEMPR12[6] ), .B(\Z\R_DATA_TEMPR13[6] ), 
        .C(\Z\R_DATA_TEMPR14[6] ), .D(\Z\R_DATA_TEMPR15[6] ), .Y(
        OR4_174_Y));
    OR2 OR2_34 (.A(\Z\R_DATA_TEMPR20[63] ), .B(\Z\R_DATA_TEMPR21[63] ), 
        .Y(OR2_34_Y));
    OR4 OR4_485 (.A(\Z\R_DATA_TEMPR8[20] ), .B(\Z\R_DATA_TEMPR9[20] ), 
        .C(\Z\R_DATA_TEMPR10[20] ), .D(\Z\R_DATA_TEMPR11[20] ), .Y(
        OR4_485_Y));
    OR4 OR4_568 (.A(\Z\R_DATA_TEMPR4[0] ), .B(\Z\R_DATA_TEMPR5[0] ), 
        .C(\Z\R_DATA_TEMPR6[0] ), .D(\Z\R_DATA_TEMPR7[0] ), .Y(
        OR4_568_Y));
    OR4 OR4_56 (.A(\Z\R_DATA_TEMPR16[4] ), .B(\Z\R_DATA_TEMPR17[4] ), 
        .C(\Z\R_DATA_TEMPR18[4] ), .D(\Z\R_DATA_TEMPR19[4] ), .Y(
        OR4_56_Y));
    OR4 OR4_532 (.A(\Z\R_DATA_TEMPR24[58] ), .B(\Z\R_DATA_TEMPR25[58] )
        , .C(\Z\R_DATA_TEMPR26[58] ), .D(\Z\R_DATA_TEMPR27[58] ), .Y(
        OR4_532_Y));
    OR4 OR4_390 (.A(\Z\R_DATA_TEMPR16[66] ), .B(\Z\R_DATA_TEMPR17[66] )
        , .C(\Z\R_DATA_TEMPR18[66] ), .D(\Z\R_DATA_TEMPR19[66] ), .Y(
        OR4_390_Y));
    OR2 OR2_55 (.A(\Z\R_DATA_TEMPR20[19] ), .B(\Z\R_DATA_TEMPR21[19] ), 
        .Y(OR2_55_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[2]  (.A(CFG2_1_Y), .B(
        R_ADDR_c[13]), .C(R_EN_c), .Y(\Z\BLKY2[2] ));
    OR4 OR4_701 (.A(\Z\R_DATA_TEMPR24[35] ), .B(\Z\R_DATA_TEMPR25[35] )
        , .C(\Z\R_DATA_TEMPR26[35] ), .D(\Z\R_DATA_TEMPR27[35] ), .Y(
        OR4_701_Y));
    OR4 \OR4_R_DATA[2]  (.A(OR4_392_Y), .B(OR4_358_Y), .C(OR4_499_Y), 
        .D(OR4_551_Y), .Y(R_DATA_c[2]));
    OR4 OR4_521 (.A(OR4_389_Y), .B(OR2_75_Y), .C(
        \Z\R_DATA_TEMPR22[53] ), .D(\Z\R_DATA_TEMPR23[53] ), .Y(
        OR4_521_Y));
    OR4 OR4_152 (.A(\Z\R_DATA_TEMPR12[54] ), .B(\Z\R_DATA_TEMPR13[54] )
        , .C(\Z\R_DATA_TEMPR14[54] ), .D(\Z\R_DATA_TEMPR15[54] ), .Y(
        OR4_152_Y));
    OR4 OR4_466 (.A(\Z\R_DATA_TEMPR8[23] ), .B(\Z\R_DATA_TEMPR9[23] ), 
        .C(\Z\R_DATA_TEMPR10[23] ), .D(\Z\R_DATA_TEMPR11[23] ), .Y(
        OR4_466_Y));
    OR4 OR4_39 (.A(\Z\R_DATA_TEMPR24[74] ), .B(\Z\R_DATA_TEMPR25[74] ), 
        .C(\Z\R_DATA_TEMPR26[74] ), .D(\Z\R_DATA_TEMPR27[74] ), .Y(
        OR4_39_Y));
    OR4 OR4_534 (.A(OR4_475_Y), .B(OR4_317_Y), .C(OR4_485_Y), .D(
        OR4_82_Y), .Y(OR4_534_Y));
    OR4 OR4_506 (.A(\Z\R_DATA_TEMPR0[70] ), .B(\Z\R_DATA_TEMPR1[70] ), 
        .C(\Z\R_DATA_TEMPR2[70] ), .D(\Z\R_DATA_TEMPR3[70] ), .Y(
        OR4_506_Y));
    OR4 OR4_211 (.A(\Z\R_DATA_TEMPR16[7] ), .B(\Z\R_DATA_TEMPR17[7] ), 
        .C(\Z\R_DATA_TEMPR18[7] ), .D(\Z\R_DATA_TEMPR19[7] ), .Y(
        OR4_211_Y));
    OR4 OR4_484 (.A(\Z\R_DATA_TEMPR0[57] ), .B(\Z\R_DATA_TEMPR1[57] ), 
        .C(\Z\R_DATA_TEMPR2[57] ), .D(\Z\R_DATA_TEMPR3[57] ), .Y(
        OR4_484_Y));
    OR2 OR2_9 (.A(\Z\R_DATA_TEMPR20[26] ), .B(\Z\R_DATA_TEMPR21[26] ), 
        .Y(OR2_9_Y));
    OR4 OR4_576 (.A(\Z\R_DATA_TEMPR4[62] ), .B(\Z\R_DATA_TEMPR5[62] ), 
        .C(\Z\R_DATA_TEMPR6[62] ), .D(\Z\R_DATA_TEMPR7[62] ), .Y(
        OR4_576_Y));
    OR4 OR4_362 (.A(OR4_100_Y), .B(OR4_149_Y), .C(OR4_387_Y), .D(
        OR4_143_Y), .Y(OR4_362_Y));
    OR4 OR4_222 (.A(\Z\R_DATA_TEMPR16[18] ), .B(\Z\R_DATA_TEMPR17[18] )
        , .C(\Z\R_DATA_TEMPR18[18] ), .D(\Z\R_DATA_TEMPR19[18] ), .Y(
        OR4_222_Y));
    OR4 OR4_145 (.A(\Z\R_DATA_TEMPR12[10] ), .B(\Z\R_DATA_TEMPR13[10] )
        , .C(\Z\R_DATA_TEMPR14[10] ), .D(\Z\R_DATA_TEMPR15[10] ), .Y(
        OR4_145_Y));
    OR4 OR4_386 (.A(\Z\R_DATA_TEMPR16[19] ), .B(\Z\R_DATA_TEMPR17[19] )
        , .C(\Z\R_DATA_TEMPR18[19] ), .D(\Z\R_DATA_TEMPR19[19] ), .Y(
        OR4_386_Y));
    OR4 OR4_16 (.A(\Z\R_DATA_TEMPR12[1] ), .B(\Z\R_DATA_TEMPR13[1] ), 
        .C(\Z\R_DATA_TEMPR14[1] ), .D(\Z\R_DATA_TEMPR15[1] ), .Y(
        OR4_16_Y));
    OR4 OR4_447 (.A(\Z\R_DATA_TEMPR28[71] ), .B(\Z\R_DATA_TEMPR29[71] )
        , .C(\Z\R_DATA_TEMPR30[71] ), .D(\Z\R_DATA_TEMPR31[71] ), .Y(
        OR4_447_Y));
    OR4 OR4_259 (.A(\Z\R_DATA_TEMPR8[34] ), .B(\Z\R_DATA_TEMPR9[34] ), 
        .C(\Z\R_DATA_TEMPR10[34] ), .D(\Z\R_DATA_TEMPR11[34] ), .Y(
        OR4_259_Y));
    OR4 OR4_4 (.A(\Z\R_DATA_TEMPR24[24] ), .B(\Z\R_DATA_TEMPR25[24] ), 
        .C(\Z\R_DATA_TEMPR26[24] ), .D(\Z\R_DATA_TEMPR27[24] ), .Y(
        OR4_4_Y));
    OR4 OR4_331 (.A(\Z\R_DATA_TEMPR16[27] ), .B(\Z\R_DATA_TEMPR17[27] )
        , .C(\Z\R_DATA_TEMPR18[27] ), .D(\Z\R_DATA_TEMPR19[27] ), .Y(
        OR4_331_Y));
    OR4 OR4_512 (.A(\Z\R_DATA_TEMPR12[17] ), .B(\Z\R_DATA_TEMPR13[17] )
        , .C(\Z\R_DATA_TEMPR14[17] ), .D(\Z\R_DATA_TEMPR15[17] ), .Y(
        OR4_512_Y));
    OR4 OR4_320 (.A(\Z\R_DATA_TEMPR28[15] ), .B(\Z\R_DATA_TEMPR29[15] )
        , .C(\Z\R_DATA_TEMPR30[15] ), .D(\Z\R_DATA_TEMPR31[15] ), .Y(
        OR4_320_Y));
    OR4 OR4_430 (.A(\Z\R_DATA_TEMPR24[44] ), .B(\Z\R_DATA_TEMPR25[44] )
        , .C(\Z\R_DATA_TEMPR26[44] ), .D(\Z\R_DATA_TEMPR27[44] ), .Y(
        OR4_430_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%7%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0 (
        .A_DOUT({\Z\R_DATA_TEMPR7[39] , \Z\R_DATA_TEMPR7[38] , 
        \Z\R_DATA_TEMPR7[37] , \Z\R_DATA_TEMPR7[36] , 
        \Z\R_DATA_TEMPR7[35] , \Z\R_DATA_TEMPR7[34] , 
        \Z\R_DATA_TEMPR7[33] , \Z\R_DATA_TEMPR7[32] , 
        \Z\R_DATA_TEMPR7[31] , \Z\R_DATA_TEMPR7[30] , 
        \Z\R_DATA_TEMPR7[29] , \Z\R_DATA_TEMPR7[28] , 
        \Z\R_DATA_TEMPR7[27] , \Z\R_DATA_TEMPR7[26] , 
        \Z\R_DATA_TEMPR7[25] , \Z\R_DATA_TEMPR7[24] , 
        \Z\R_DATA_TEMPR7[23] , \Z\R_DATA_TEMPR7[22] , 
        \Z\R_DATA_TEMPR7[21] , \Z\R_DATA_TEMPR7[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR7[19] , \Z\R_DATA_TEMPR7[18] , 
        \Z\R_DATA_TEMPR7[17] , \Z\R_DATA_TEMPR7[16] , 
        \Z\R_DATA_TEMPR7[15] , \Z\R_DATA_TEMPR7[14] , 
        \Z\R_DATA_TEMPR7[13] , \Z\R_DATA_TEMPR7[12] , 
        \Z\R_DATA_TEMPR7[11] , \Z\R_DATA_TEMPR7[10] , 
        \Z\R_DATA_TEMPR7[9] , \Z\R_DATA_TEMPR7[8] , 
        \Z\R_DATA_TEMPR7[7] , \Z\R_DATA_TEMPR7[6] , 
        \Z\R_DATA_TEMPR7[5] , \Z\R_DATA_TEMPR7[4] , 
        \Z\R_DATA_TEMPR7[3] , \Z\R_DATA_TEMPR7[2] , 
        \Z\R_DATA_TEMPR7[1] , \Z\R_DATA_TEMPR7[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[7][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[1] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[1] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[14]  (.A(OR4_686_Y), .B(OR4_428_Y), .C(OR4_60_Y), 
        .D(OR4_380_Y), .Y(R_DATA_c[14]));
    OR4 OR4_595 (.A(\Z\R_DATA_TEMPR28[79] ), .B(\Z\R_DATA_TEMPR29[79] )
        , .C(\Z\R_DATA_TEMPR30[79] ), .D(\Z\R_DATA_TEMPR31[79] ), .Y(
        OR4_595_Y));
    OR4 OR4_245 (.A(\Z\R_DATA_TEMPR0[56] ), .B(\Z\R_DATA_TEMPR1[56] ), 
        .C(\Z\R_DATA_TEMPR2[56] ), .D(\Z\R_DATA_TEMPR3[56] ), .Y(
        OR4_245_Y));
    OR4 OR4_508 (.A(\Z\R_DATA_TEMPR8[12] ), .B(\Z\R_DATA_TEMPR9[12] ), 
        .C(\Z\R_DATA_TEMPR10[12] ), .D(\Z\R_DATA_TEMPR11[12] ), .Y(
        OR4_508_Y));
    OR4 OR4_50 (.A(\Z\R_DATA_TEMPR4[35] ), .B(\Z\R_DATA_TEMPR5[35] ), 
        .C(\Z\R_DATA_TEMPR6[35] ), .D(\Z\R_DATA_TEMPR7[35] ), .Y(
        OR4_50_Y));
    OR4 OR4_514 (.A(\Z\R_DATA_TEMPR12[53] ), .B(\Z\R_DATA_TEMPR13[53] )
        , .C(\Z\R_DATA_TEMPR14[53] ), .D(\Z\R_DATA_TEMPR15[53] ), .Y(
        OR4_514_Y));
    OR4 OR4_578 (.A(\Z\R_DATA_TEMPR24[60] ), .B(\Z\R_DATA_TEMPR25[60] )
        , .C(\Z\R_DATA_TEMPR26[60] ), .D(\Z\R_DATA_TEMPR27[60] ), .Y(
        OR4_578_Y));
    OR4 OR4_693 (.A(\Z\R_DATA_TEMPR8[33] ), .B(\Z\R_DATA_TEMPR9[33] ), 
        .C(\Z\R_DATA_TEMPR10[33] ), .D(\Z\R_DATA_TEMPR11[33] ), .Y(
        OR4_693_Y));
    OR4 OR4_57 (.A(\Z\R_DATA_TEMPR16[23] ), .B(\Z\R_DATA_TEMPR17[23] ), 
        .C(\Z\R_DATA_TEMPR18[23] ), .D(\Z\R_DATA_TEMPR19[23] ), .Y(
        OR4_57_Y));
    OR4 OR4_32 (.A(\Z\R_DATA_TEMPR28[44] ), .B(\Z\R_DATA_TEMPR29[44] ), 
        .C(\Z\R_DATA_TEMPR30[44] ), .D(\Z\R_DATA_TEMPR31[44] ), .Y(
        OR4_32_Y));
    OR4 OR4_260 (.A(\Z\R_DATA_TEMPR12[13] ), .B(\Z\R_DATA_TEMPR13[13] )
        , .C(\Z\R_DATA_TEMPR14[13] ), .D(\Z\R_DATA_TEMPR15[13] ), .Y(
        OR4_260_Y));
    OR4 OR4_567 (.A(\Z\R_DATA_TEMPR24[32] ), .B(\Z\R_DATA_TEMPR25[32] )
        , .C(\Z\R_DATA_TEMPR26[32] ), .D(\Z\R_DATA_TEMPR27[32] ), .Y(
        OR4_567_Y));
    OR4 OR4_406 (.A(\Z\R_DATA_TEMPR16[50] ), .B(\Z\R_DATA_TEMPR17[50] )
        , .C(\Z\R_DATA_TEMPR18[50] ), .D(\Z\R_DATA_TEMPR19[50] ), .Y(
        OR4_406_Y));
    OR4 OR4_443 (.A(\Z\R_DATA_TEMPR12[7] ), .B(\Z\R_DATA_TEMPR13[7] ), 
        .C(\Z\R_DATA_TEMPR14[7] ), .D(\Z\R_DATA_TEMPR15[7] ), .Y(
        OR4_443_Y));
    OR4 OR4_669 (.A(OR4_200_Y), .B(OR4_308_Y), .C(OR4_307_Y), .D(
        OR4_423_Y), .Y(OR4_669_Y));
    OR4 OR4_641 (.A(\Z\R_DATA_TEMPR24[48] ), .B(\Z\R_DATA_TEMPR25[48] )
        , .C(\Z\R_DATA_TEMPR26[48] ), .D(\Z\R_DATA_TEMPR27[48] ), .Y(
        OR4_641_Y));
    OR4 OR4_476 (.A(OR4_165_Y), .B(OR2_64_Y), .C(
        \Z\R_DATA_TEMPR22[72] ), .D(\Z\R_DATA_TEMPR23[72] ), .Y(
        OR4_476_Y));
    OR4 OR4_311 (.A(\Z\R_DATA_TEMPR12[30] ), .B(\Z\R_DATA_TEMPR13[30] )
        , .C(\Z\R_DATA_TEMPR14[30] ), .D(\Z\R_DATA_TEMPR15[30] ), .Y(
        OR4_311_Y));
    OR4 OR4_184 (.A(\Z\R_DATA_TEMPR0[63] ), .B(\Z\R_DATA_TEMPR1[63] ), 
        .C(\Z\R_DATA_TEMPR2[63] ), .D(\Z\R_DATA_TEMPR3[63] ), .Y(
        OR4_184_Y));
    OR4 OR4_248 (.A(\Z\R_DATA_TEMPR24[78] ), .B(\Z\R_DATA_TEMPR25[78] )
        , .C(\Z\R_DATA_TEMPR26[78] ), .D(\Z\R_DATA_TEMPR27[78] ), .Y(
        OR4_248_Y));
    OR4 OR4_302 (.A(\Z\R_DATA_TEMPR24[36] ), .B(\Z\R_DATA_TEMPR25[36] )
        , .C(\Z\R_DATA_TEMPR26[36] ), .D(\Z\R_DATA_TEMPR27[36] ), .Y(
        OR4_302_Y));
    OR4 OR4_266 (.A(OR4_113_Y), .B(OR2_76_Y), .C(
        \Z\R_DATA_TEMPR22[13] ), .D(\Z\R_DATA_TEMPR23[13] ), .Y(
        OR4_266_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%8%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C1 (
        .A_DOUT({\Z\R_DATA_TEMPR8[79] , \Z\R_DATA_TEMPR8[78] , 
        \Z\R_DATA_TEMPR8[77] , \Z\R_DATA_TEMPR8[76] , 
        \Z\R_DATA_TEMPR8[75] , \Z\R_DATA_TEMPR8[74] , 
        \Z\R_DATA_TEMPR8[73] , \Z\R_DATA_TEMPR8[72] , 
        \Z\R_DATA_TEMPR8[71] , \Z\R_DATA_TEMPR8[70] , 
        \Z\R_DATA_TEMPR8[69] , \Z\R_DATA_TEMPR8[68] , 
        \Z\R_DATA_TEMPR8[67] , \Z\R_DATA_TEMPR8[66] , 
        \Z\R_DATA_TEMPR8[65] , \Z\R_DATA_TEMPR8[64] , 
        \Z\R_DATA_TEMPR8[63] , \Z\R_DATA_TEMPR8[62] , 
        \Z\R_DATA_TEMPR8[61] , \Z\R_DATA_TEMPR8[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR8[59] , \Z\R_DATA_TEMPR8[58] , 
        \Z\R_DATA_TEMPR8[57] , \Z\R_DATA_TEMPR8[56] , 
        \Z\R_DATA_TEMPR8[55] , \Z\R_DATA_TEMPR8[54] , 
        \Z\R_DATA_TEMPR8[53] , \Z\R_DATA_TEMPR8[52] , 
        \Z\R_DATA_TEMPR8[51] , \Z\R_DATA_TEMPR8[50] , 
        \Z\R_DATA_TEMPR8[49] , \Z\R_DATA_TEMPR8[48] , 
        \Z\R_DATA_TEMPR8[47] , \Z\R_DATA_TEMPR8[46] , 
        \Z\R_DATA_TEMPR8[45] , \Z\R_DATA_TEMPR8[44] , 
        \Z\R_DATA_TEMPR8[43] , \Z\R_DATA_TEMPR8[42] , 
        \Z\R_DATA_TEMPR8[41] , \Z\R_DATA_TEMPR8[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[8][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[2] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[2] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_76 (.A(\Z\R_DATA_TEMPR28[10] ), .B(\Z\R_DATA_TEMPR29[10] ), 
        .C(\Z\R_DATA_TEMPR30[10] ), .D(\Z\R_DATA_TEMPR31[10] ), .Y(
        OR4_76_Y));
    OR4 OR4_410 (.A(\Z\R_DATA_TEMPR4[49] ), .B(\Z\R_DATA_TEMPR5[49] ), 
        .C(\Z\R_DATA_TEMPR6[49] ), .D(\Z\R_DATA_TEMPR7[49] ), .Y(
        OR4_410_Y));
    OR4 OR4_25 (.A(\Z\R_DATA_TEMPR28[51] ), .B(\Z\R_DATA_TEMPR29[51] ), 
        .C(\Z\R_DATA_TEMPR30[51] ), .D(\Z\R_DATA_TEMPR31[51] ), .Y(
        OR4_25_Y));
    OR4 OR4_10 (.A(\Z\R_DATA_TEMPR24[40] ), .B(\Z\R_DATA_TEMPR25[40] ), 
        .C(\Z\R_DATA_TEMPR26[40] ), .D(\Z\R_DATA_TEMPR27[40] ), .Y(
        OR4_10_Y));
    OR4 OR4_339 (.A(\Z\R_DATA_TEMPR24[22] ), .B(\Z\R_DATA_TEMPR25[22] )
        , .C(\Z\R_DATA_TEMPR26[22] ), .D(\Z\R_DATA_TEMPR27[22] ), .Y(
        OR4_339_Y));
    OR4 OR4_193 (.A(OR4_394_Y), .B(OR2_63_Y), .C(
        \Z\R_DATA_TEMPR22[61] ), .D(\Z\R_DATA_TEMPR23[61] ), .Y(
        OR4_193_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[4]  (.A(CFG2_4_Y), .B(
        W_ADDR_c[13]), .C(W_EN_c), .Y(\Z\BLKX2[4] ));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%4%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C1 (
        .A_DOUT({\Z\R_DATA_TEMPR4[79] , \Z\R_DATA_TEMPR4[78] , 
        \Z\R_DATA_TEMPR4[77] , \Z\R_DATA_TEMPR4[76] , 
        \Z\R_DATA_TEMPR4[75] , \Z\R_DATA_TEMPR4[74] , 
        \Z\R_DATA_TEMPR4[73] , \Z\R_DATA_TEMPR4[72] , 
        \Z\R_DATA_TEMPR4[71] , \Z\R_DATA_TEMPR4[70] , 
        \Z\R_DATA_TEMPR4[69] , \Z\R_DATA_TEMPR4[68] , 
        \Z\R_DATA_TEMPR4[67] , \Z\R_DATA_TEMPR4[66] , 
        \Z\R_DATA_TEMPR4[65] , \Z\R_DATA_TEMPR4[64] , 
        \Z\R_DATA_TEMPR4[63] , \Z\R_DATA_TEMPR4[62] , 
        \Z\R_DATA_TEMPR4[61] , \Z\R_DATA_TEMPR4[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR4[59] , \Z\R_DATA_TEMPR4[58] , 
        \Z\R_DATA_TEMPR4[57] , \Z\R_DATA_TEMPR4[56] , 
        \Z\R_DATA_TEMPR4[55] , \Z\R_DATA_TEMPR4[54] , 
        \Z\R_DATA_TEMPR4[53] , \Z\R_DATA_TEMPR4[52] , 
        \Z\R_DATA_TEMPR4[51] , \Z\R_DATA_TEMPR4[50] , 
        \Z\R_DATA_TEMPR4[49] , \Z\R_DATA_TEMPR4[48] , 
        \Z\R_DATA_TEMPR4[47] , \Z\R_DATA_TEMPR4[46] , 
        \Z\R_DATA_TEMPR4[45] , \Z\R_DATA_TEMPR4[44] , 
        \Z\R_DATA_TEMPR4[43] , \Z\R_DATA_TEMPR4[42] , 
        \Z\R_DATA_TEMPR4[41] , \Z\R_DATA_TEMPR4[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[4][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[1] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[1] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_372 (.A(\Z\R_DATA_TEMPR24[72] ), .B(\Z\R_DATA_TEMPR25[72] )
        , .C(\Z\R_DATA_TEMPR26[72] ), .D(\Z\R_DATA_TEMPR27[72] ), .Y(
        OR4_372_Y));
    OR4 \OR4_R_DATA[44]  (.A(OR4_335_Y), .B(OR4_84_Y), .C(OR4_430_Y), 
        .D(OR4_32_Y), .Y(R_DATA_c[44]));
    OR4 OR4_525 (.A(\Z\R_DATA_TEMPR8[0] ), .B(\Z\R_DATA_TEMPR9[0] ), 
        .C(\Z\R_DATA_TEMPR10[0] ), .D(\Z\R_DATA_TEMPR11[0] ), .Y(
        OR4_525_Y));
    OR4 OR4_17 (.A(\Z\R_DATA_TEMPR4[56] ), .B(\Z\R_DATA_TEMPR5[56] ), 
        .C(\Z\R_DATA_TEMPR6[56] ), .D(\Z\R_DATA_TEMPR7[56] ), .Y(
        OR4_17_Y));
    OR4 OR4_664 (.A(OR4_150_Y), .B(OR2_3_Y), .C(\Z\R_DATA_TEMPR22[71] )
        , .D(\Z\R_DATA_TEMPR23[71] ), .Y(OR4_664_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%13%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C1 (
        .A_DOUT({\Z\R_DATA_TEMPR13[79] , \Z\R_DATA_TEMPR13[78] , 
        \Z\R_DATA_TEMPR13[77] , \Z\R_DATA_TEMPR13[76] , 
        \Z\R_DATA_TEMPR13[75] , \Z\R_DATA_TEMPR13[74] , 
        \Z\R_DATA_TEMPR13[73] , \Z\R_DATA_TEMPR13[72] , 
        \Z\R_DATA_TEMPR13[71] , \Z\R_DATA_TEMPR13[70] , 
        \Z\R_DATA_TEMPR13[69] , \Z\R_DATA_TEMPR13[68] , 
        \Z\R_DATA_TEMPR13[67] , \Z\R_DATA_TEMPR13[66] , 
        \Z\R_DATA_TEMPR13[65] , \Z\R_DATA_TEMPR13[64] , 
        \Z\R_DATA_TEMPR13[63] , \Z\R_DATA_TEMPR13[62] , 
        \Z\R_DATA_TEMPR13[61] , \Z\R_DATA_TEMPR13[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR13[59] , \Z\R_DATA_TEMPR13[58] , 
        \Z\R_DATA_TEMPR13[57] , \Z\R_DATA_TEMPR13[56] , 
        \Z\R_DATA_TEMPR13[55] , \Z\R_DATA_TEMPR13[54] , 
        \Z\R_DATA_TEMPR13[53] , \Z\R_DATA_TEMPR13[52] , 
        \Z\R_DATA_TEMPR13[51] , \Z\R_DATA_TEMPR13[50] , 
        \Z\R_DATA_TEMPR13[49] , \Z\R_DATA_TEMPR13[48] , 
        \Z\R_DATA_TEMPR13[47] , \Z\R_DATA_TEMPR13[46] , 
        \Z\R_DATA_TEMPR13[45] , \Z\R_DATA_TEMPR13[44] , 
        \Z\R_DATA_TEMPR13[43] , \Z\R_DATA_TEMPR13[42] , 
        \Z\R_DATA_TEMPR13[41] , \Z\R_DATA_TEMPR13[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[13][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[3] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[3] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_623 (.A(\Z\R_DATA_TEMPR0[41] ), .B(\Z\R_DATA_TEMPR1[41] ), 
        .C(\Z\R_DATA_TEMPR2[41] ), .D(\Z\R_DATA_TEMPR3[41] ), .Y(
        OR4_623_Y));
    OR4 OR4_586 (.A(\Z\R_DATA_TEMPR8[61] ), .B(\Z\R_DATA_TEMPR9[61] ), 
        .C(\Z\R_DATA_TEMPR10[61] ), .D(\Z\R_DATA_TEMPR11[61] ), .Y(
        OR4_586_Y));
    OR4 OR4_200 (.A(\Z\R_DATA_TEMPR0[21] ), .B(\Z\R_DATA_TEMPR1[21] ), 
        .C(\Z\R_DATA_TEMPR2[21] ), .D(\Z\R_DATA_TEMPR3[21] ), .Y(
        OR4_200_Y));
    OR4 \OR4_R_DATA[64]  (.A(OR4_189_Y), .B(OR4_652_Y), .C(OR4_283_Y), 
        .D(OR4_598_Y), .Y(R_DATA_c[64]));
    OR4 OR4_507 (.A(\Z\R_DATA_TEMPR4[73] ), .B(\Z\R_DATA_TEMPR5[73] ), 
        .C(\Z\R_DATA_TEMPR6[73] ), .D(\Z\R_DATA_TEMPR7[73] ), .Y(
        OR4_507_Y));
    OR2 OR2_59 (.A(\Z\R_DATA_TEMPR20[46] ), .B(\Z\R_DATA_TEMPR21[46] ), 
        .Y(OR2_59_Y));
    OR4 OR4_270 (.A(\Z\R_DATA_TEMPR12[44] ), .B(\Z\R_DATA_TEMPR13[44] )
        , .C(\Z\R_DATA_TEMPR14[44] ), .D(\Z\R_DATA_TEMPR15[44] ), .Y(
        OR4_270_Y));
    OR4 OR4_577 (.A(\Z\R_DATA_TEMPR28[43] ), .B(\Z\R_DATA_TEMPR29[43] )
        , .C(\Z\R_DATA_TEMPR30[43] ), .D(\Z\R_DATA_TEMPR31[43] ), .Y(
        OR4_577_Y));
    OR4 OR4_541 (.A(\Z\R_DATA_TEMPR4[13] ), .B(\Z\R_DATA_TEMPR5[13] ), 
        .C(\Z\R_DATA_TEMPR6[13] ), .D(\Z\R_DATA_TEMPR7[13] ), .Y(
        OR4_541_Y));
    OR4 OR4_319 (.A(\Z\R_DATA_TEMPR16[29] ), .B(\Z\R_DATA_TEMPR17[29] )
        , .C(\Z\R_DATA_TEMPR18[29] ), .D(\Z\R_DATA_TEMPR19[29] ), .Y(
        OR4_319_Y));
    OR4 OR4_192 (.A(\Z\R_DATA_TEMPR12[56] ), .B(\Z\R_DATA_TEMPR13[56] )
        , .C(\Z\R_DATA_TEMPR14[56] ), .D(\Z\R_DATA_TEMPR15[56] ), .Y(
        OR4_192_Y));
    OR4 OR4_609 (.A(\Z\R_DATA_TEMPR12[48] ), .B(\Z\R_DATA_TEMPR13[48] )
        , .C(\Z\R_DATA_TEMPR14[48] ), .D(\Z\R_DATA_TEMPR15[48] ), .Y(
        OR4_609_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%28%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C1 (
        .A_DOUT({\Z\R_DATA_TEMPR28[79] , \Z\R_DATA_TEMPR28[78] , 
        \Z\R_DATA_TEMPR28[77] , \Z\R_DATA_TEMPR28[76] , 
        \Z\R_DATA_TEMPR28[75] , \Z\R_DATA_TEMPR28[74] , 
        \Z\R_DATA_TEMPR28[73] , \Z\R_DATA_TEMPR28[72] , 
        \Z\R_DATA_TEMPR28[71] , \Z\R_DATA_TEMPR28[70] , 
        \Z\R_DATA_TEMPR28[69] , \Z\R_DATA_TEMPR28[68] , 
        \Z\R_DATA_TEMPR28[67] , \Z\R_DATA_TEMPR28[66] , 
        \Z\R_DATA_TEMPR28[65] , \Z\R_DATA_TEMPR28[64] , 
        \Z\R_DATA_TEMPR28[63] , \Z\R_DATA_TEMPR28[62] , 
        \Z\R_DATA_TEMPR28[61] , \Z\R_DATA_TEMPR28[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR28[59] , \Z\R_DATA_TEMPR28[58] , 
        \Z\R_DATA_TEMPR28[57] , \Z\R_DATA_TEMPR28[56] , 
        \Z\R_DATA_TEMPR28[55] , \Z\R_DATA_TEMPR28[54] , 
        \Z\R_DATA_TEMPR28[53] , \Z\R_DATA_TEMPR28[52] , 
        \Z\R_DATA_TEMPR28[51] , \Z\R_DATA_TEMPR28[50] , 
        \Z\R_DATA_TEMPR28[49] , \Z\R_DATA_TEMPR28[48] , 
        \Z\R_DATA_TEMPR28[47] , \Z\R_DATA_TEMPR28[46] , 
        \Z\R_DATA_TEMPR28[45] , \Z\R_DATA_TEMPR28[44] , 
        \Z\R_DATA_TEMPR28[43] , \Z\R_DATA_TEMPR28[42] , 
        \Z\R_DATA_TEMPR28[41] , \Z\R_DATA_TEMPR28[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[28][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[7] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[7] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_123 (.A(\Z\R_DATA_TEMPR0[25] ), .B(\Z\R_DATA_TEMPR1[25] ), 
        .C(\Z\R_DATA_TEMPR2[25] ), .D(\Z\R_DATA_TEMPR3[25] ), .Y(
        OR4_123_Y));
    OR4 OR4_679 (.A(\Z\R_DATA_TEMPR0[13] ), .B(\Z\R_DATA_TEMPR1[13] ), 
        .C(\Z\R_DATA_TEMPR2[13] ), .D(\Z\R_DATA_TEMPR3[13] ), .Y(
        OR4_679_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%14%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0 (
        .A_DOUT({\Z\R_DATA_TEMPR14[39] , \Z\R_DATA_TEMPR14[38] , 
        \Z\R_DATA_TEMPR14[37] , \Z\R_DATA_TEMPR14[36] , 
        \Z\R_DATA_TEMPR14[35] , \Z\R_DATA_TEMPR14[34] , 
        \Z\R_DATA_TEMPR14[33] , \Z\R_DATA_TEMPR14[32] , 
        \Z\R_DATA_TEMPR14[31] , \Z\R_DATA_TEMPR14[30] , 
        \Z\R_DATA_TEMPR14[29] , \Z\R_DATA_TEMPR14[28] , 
        \Z\R_DATA_TEMPR14[27] , \Z\R_DATA_TEMPR14[26] , 
        \Z\R_DATA_TEMPR14[25] , \Z\R_DATA_TEMPR14[24] , 
        \Z\R_DATA_TEMPR14[23] , \Z\R_DATA_TEMPR14[22] , 
        \Z\R_DATA_TEMPR14[21] , \Z\R_DATA_TEMPR14[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR14[19] , \Z\R_DATA_TEMPR14[18] , 
        \Z\R_DATA_TEMPR14[17] , \Z\R_DATA_TEMPR14[16] , 
        \Z\R_DATA_TEMPR14[15] , \Z\R_DATA_TEMPR14[14] , 
        \Z\R_DATA_TEMPR14[13] , \Z\R_DATA_TEMPR14[12] , 
        \Z\R_DATA_TEMPR14[11] , \Z\R_DATA_TEMPR14[10] , 
        \Z\R_DATA_TEMPR14[9] , \Z\R_DATA_TEMPR14[8] , 
        \Z\R_DATA_TEMPR14[7] , \Z\R_DATA_TEMPR14[6] , 
        \Z\R_DATA_TEMPR14[5] , \Z\R_DATA_TEMPR14[4] , 
        \Z\R_DATA_TEMPR14[3] , \Z\R_DATA_TEMPR14[2] , 
        \Z\R_DATA_TEMPR14[1] , \Z\R_DATA_TEMPR14[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[14][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[3] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[3] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_206 (.A(OR4_57_Y), .B(OR2_24_Y), .C(\Z\R_DATA_TEMPR22[23] )
        , .D(\Z\R_DATA_TEMPR23[23] ), .Y(OR4_206_Y));
    OR4 OR4_533 (.A(\Z\R_DATA_TEMPR8[7] ), .B(\Z\R_DATA_TEMPR9[7] ), 
        .C(\Z\R_DATA_TEMPR10[7] ), .D(\Z\R_DATA_TEMPR11[7] ), .Y(
        OR4_533_Y));
    OR4 OR4_70 (.A(\Z\R_DATA_TEMPR24[55] ), .B(\Z\R_DATA_TEMPR25[55] ), 
        .C(\Z\R_DATA_TEMPR26[55] ), .D(\Z\R_DATA_TEMPR27[55] ), .Y(
        OR4_70_Y));
    CFG2 #( .INIT(4'h2) )  CFG2_1 (.A(R_ADDR_c[12]), .B(R_ADDR_c[11]), 
        .Y(CFG2_1_Y));
    OR4 OR4_588 (.A(\Z\R_DATA_TEMPR4[58] ), .B(\Z\R_DATA_TEMPR5[58] ), 
        .C(\Z\R_DATA_TEMPR6[58] ), .D(\Z\R_DATA_TEMPR7[58] ), .Y(
        OR4_588_Y));
    OR4 OR4_58 (.A(\Z\R_DATA_TEMPR28[39] ), .B(\Z\R_DATA_TEMPR29[39] ), 
        .C(\Z\R_DATA_TEMPR30[39] ), .D(\Z\R_DATA_TEMPR31[39] ), .Y(
        OR4_58_Y));
    OR4 OR4_276 (.A(\Z\R_DATA_TEMPR4[54] ), .B(\Z\R_DATA_TEMPR5[54] ), 
        .C(\Z\R_DATA_TEMPR6[54] ), .D(\Z\R_DATA_TEMPR7[54] ), .Y(
        OR4_276_Y));
    OR4 OR4_77 (.A(\Z\R_DATA_TEMPR8[35] ), .B(\Z\R_DATA_TEMPR9[35] ), 
        .C(\Z\R_DATA_TEMPR10[35] ), .D(\Z\R_DATA_TEMPR11[35] ), .Y(
        OR4_77_Y));
    OR4 OR4_242 (.A(OR4_375_Y), .B(OR2_10_Y), .C(\Z\R_DATA_TEMPR22[9] )
        , .D(\Z\R_DATA_TEMPR23[9] ), .Y(OR4_242_Y));
    OR4 OR4_604 (.A(OR4_65_Y), .B(OR2_36_Y), .C(\Z\R_DATA_TEMPR22[34] )
        , .D(\Z\R_DATA_TEMPR23[34] ), .Y(OR4_604_Y));
    OR4 OR4_299 (.A(\Z\R_DATA_TEMPR28[60] ), .B(\Z\R_DATA_TEMPR29[60] )
        , .C(\Z\R_DATA_TEMPR30[60] ), .D(\Z\R_DATA_TEMPR31[60] ), .Y(
        OR4_299_Y));
    OR4 OR4_674 (.A(\Z\R_DATA_TEMPR24[71] ), .B(\Z\R_DATA_TEMPR25[71] )
        , .C(\Z\R_DATA_TEMPR26[71] ), .D(\Z\R_DATA_TEMPR27[71] ), .Y(
        OR4_674_Y));
    OR4 OR4_455 (.A(\Z\R_DATA_TEMPR12[71] ), .B(\Z\R_DATA_TEMPR13[71] )
        , .C(\Z\R_DATA_TEMPR14[71] ), .D(\Z\R_DATA_TEMPR15[71] ), .Y(
        OR4_455_Y));
    OR4 OR4_486 (.A(\Z\R_DATA_TEMPR8[72] ), .B(\Z\R_DATA_TEMPR9[72] ), 
        .C(\Z\R_DATA_TEMPR10[72] ), .D(\Z\R_DATA_TEMPR11[72] ), .Y(
        OR4_486_Y));
    OR4 \OR4_R_DATA[5]  (.A(OR4_107_Y), .B(OR4_688_Y), .C(OR4_457_Y), 
        .D(OR4_601_Y), .Y(R_DATA_c[5]));
    OR4 OR4_340 (.A(\Z\R_DATA_TEMPR16[36] ), .B(\Z\R_DATA_TEMPR17[36] )
        , .C(\Z\R_DATA_TEMPR18[36] ), .D(\Z\R_DATA_TEMPR19[36] ), .Y(
        OR4_340_Y));
    OR2 OR2_52 (.A(\Z\R_DATA_TEMPR20[28] ), .B(\Z\R_DATA_TEMPR21[28] ), 
        .Y(OR2_52_Y));
    OR4 OR4_719 (.A(\Z\R_DATA_TEMPR8[49] ), .B(\Z\R_DATA_TEMPR9[49] ), 
        .C(\Z\R_DATA_TEMPR10[49] ), .D(\Z\R_DATA_TEMPR11[49] ), .Y(
        OR4_719_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%26%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C1 (
        .A_DOUT({\Z\R_DATA_TEMPR26[79] , \Z\R_DATA_TEMPR26[78] , 
        \Z\R_DATA_TEMPR26[77] , \Z\R_DATA_TEMPR26[76] , 
        \Z\R_DATA_TEMPR26[75] , \Z\R_DATA_TEMPR26[74] , 
        \Z\R_DATA_TEMPR26[73] , \Z\R_DATA_TEMPR26[72] , 
        \Z\R_DATA_TEMPR26[71] , \Z\R_DATA_TEMPR26[70] , 
        \Z\R_DATA_TEMPR26[69] , \Z\R_DATA_TEMPR26[68] , 
        \Z\R_DATA_TEMPR26[67] , \Z\R_DATA_TEMPR26[66] , 
        \Z\R_DATA_TEMPR26[65] , \Z\R_DATA_TEMPR26[64] , 
        \Z\R_DATA_TEMPR26[63] , \Z\R_DATA_TEMPR26[62] , 
        \Z\R_DATA_TEMPR26[61] , \Z\R_DATA_TEMPR26[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR26[59] , \Z\R_DATA_TEMPR26[58] , 
        \Z\R_DATA_TEMPR26[57] , \Z\R_DATA_TEMPR26[56] , 
        \Z\R_DATA_TEMPR26[55] , \Z\R_DATA_TEMPR26[54] , 
        \Z\R_DATA_TEMPR26[53] , \Z\R_DATA_TEMPR26[52] , 
        \Z\R_DATA_TEMPR26[51] , \Z\R_DATA_TEMPR26[50] , 
        \Z\R_DATA_TEMPR26[49] , \Z\R_DATA_TEMPR26[48] , 
        \Z\R_DATA_TEMPR26[47] , \Z\R_DATA_TEMPR26[46] , 
        \Z\R_DATA_TEMPR26[45] , \Z\R_DATA_TEMPR26[44] , 
        \Z\R_DATA_TEMPR26[43] , \Z\R_DATA_TEMPR26[42] , 
        \Z\R_DATA_TEMPR26[41] , \Z\R_DATA_TEMPR26[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[26][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[6] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[6] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[11]  (.A(OR4_2_Y), .B(OR4_691_Y), .C(OR4_706_Y), 
        .D(OR4_481_Y), .Y(R_DATA_c[11]));
    OR4 OR4_122 (.A(OR4_14_Y), .B(OR4_166_Y), .C(OR4_259_Y), .D(
        OR4_47_Y), .Y(OR4_122_Y));
    OR4 OR4_382 (.A(\Z\R_DATA_TEMPR4[10] ), .B(\Z\R_DATA_TEMPR5[10] ), 
        .C(\Z\R_DATA_TEMPR6[10] ), .D(\Z\R_DATA_TEMPR7[10] ), .Y(
        OR4_382_Y));
    OR4 \OR4_R_DATA[9]  (.A(OR4_90_Y), .B(OR4_242_Y), .C(OR4_417_Y), 
        .D(OR4_560_Y), .Y(R_DATA_c[9]));
    OR4 OR4_18 (.A(\Z\R_DATA_TEMPR28[22] ), .B(\Z\R_DATA_TEMPR29[22] ), 
        .C(\Z\R_DATA_TEMPR30[22] ), .D(\Z\R_DATA_TEMPR31[22] ), .Y(
        OR4_18_Y));
    OR4 OR4_513 (.A(\Z\R_DATA_TEMPR8[70] ), .B(\Z\R_DATA_TEMPR9[70] ), 
        .C(\Z\R_DATA_TEMPR10[70] ), .D(\Z\R_DATA_TEMPR11[70] ), .Y(
        OR4_513_Y));
    OR4 OR4_34 (.A(OR4_138_Y), .B(OR2_12_Y), .C(\Z\R_DATA_TEMPR22[10] )
        , .D(\Z\R_DATA_TEMPR23[10] ), .Y(OR4_34_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%0%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0 (
        .A_DOUT({\Z\R_DATA_TEMPR0[39] , \Z\R_DATA_TEMPR0[38] , 
        \Z\R_DATA_TEMPR0[37] , \Z\R_DATA_TEMPR0[36] , 
        \Z\R_DATA_TEMPR0[35] , \Z\R_DATA_TEMPR0[34] , 
        \Z\R_DATA_TEMPR0[33] , \Z\R_DATA_TEMPR0[32] , 
        \Z\R_DATA_TEMPR0[31] , \Z\R_DATA_TEMPR0[30] , 
        \Z\R_DATA_TEMPR0[29] , \Z\R_DATA_TEMPR0[28] , 
        \Z\R_DATA_TEMPR0[27] , \Z\R_DATA_TEMPR0[26] , 
        \Z\R_DATA_TEMPR0[25] , \Z\R_DATA_TEMPR0[24] , 
        \Z\R_DATA_TEMPR0[23] , \Z\R_DATA_TEMPR0[22] , 
        \Z\R_DATA_TEMPR0[21] , \Z\R_DATA_TEMPR0[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR0[19] , \Z\R_DATA_TEMPR0[18] , 
        \Z\R_DATA_TEMPR0[17] , \Z\R_DATA_TEMPR0[16] , 
        \Z\R_DATA_TEMPR0[15] , \Z\R_DATA_TEMPR0[14] , 
        \Z\R_DATA_TEMPR0[13] , \Z\R_DATA_TEMPR0[12] , 
        \Z\R_DATA_TEMPR0[11] , \Z\R_DATA_TEMPR0[10] , 
        \Z\R_DATA_TEMPR0[9] , \Z\R_DATA_TEMPR0[8] , 
        \Z\R_DATA_TEMPR0[7] , \Z\R_DATA_TEMPR0[6] , 
        \Z\R_DATA_TEMPR0[5] , \Z\R_DATA_TEMPR0[4] , 
        \Z\R_DATA_TEMPR0[3] , \Z\R_DATA_TEMPR0[2] , 
        \Z\R_DATA_TEMPR0[1] , \Z\R_DATA_TEMPR0[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[0][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[0] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[0] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_454 (.A(\Z\R_DATA_TEMPR28[40] ), .B(\Z\R_DATA_TEMPR29[40] )
        , .C(\Z\R_DATA_TEMPR30[40] ), .D(\Z\R_DATA_TEMPR31[40] ), .Y(
        OR4_454_Y));
    OR4 \OR4_R_DATA[35]  (.A(OR4_67_Y), .B(OR4_418_Y), .C(OR4_701_Y), 
        .D(OR4_494_Y), .Y(R_DATA_c[35]));
    OR4 \OR4_R_DATA[10]  (.A(OR4_593_Y), .B(OR4_34_Y), .C(OR4_359_Y), 
        .D(OR4_76_Y), .Y(R_DATA_c[10]));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[1]  (.A(CFG2_2_Y), .B(
        W_ADDR_c[13]), .C(W_EN_c), .Y(\Z\BLKX2[1] ));
    OR4 OR4_229 (.A(\Z\R_DATA_TEMPR0[71] ), .B(\Z\R_DATA_TEMPR1[71] ), 
        .C(\Z\R_DATA_TEMPR2[71] ), .D(\Z\R_DATA_TEMPR3[71] ), .Y(
        OR4_229_Y));
    OR4 OR4_356 (.A(\Z\R_DATA_TEMPR4[12] ), .B(\Z\R_DATA_TEMPR5[12] ), 
        .C(\Z\R_DATA_TEMPR6[12] ), .D(\Z\R_DATA_TEMPR7[12] ), .Y(
        OR4_356_Y));
    OR4 OR4_261 (.A(\Z\R_DATA_TEMPR24[51] ), .B(\Z\R_DATA_TEMPR25[51] )
        , .C(\Z\R_DATA_TEMPR26[51] ), .D(\Z\R_DATA_TEMPR27[51] ), .Y(
        OR4_261_Y));
    OR2 OR2_23 (.A(\Z\R_DATA_TEMPR20[77] ), .B(\Z\R_DATA_TEMPR21[77] ), 
        .Y(OR2_23_Y));
    OR4 OR4_29 (.A(\Z\R_DATA_TEMPR28[17] ), .B(\Z\R_DATA_TEMPR29[17] ), 
        .C(\Z\R_DATA_TEMPR30[17] ), .D(\Z\R_DATA_TEMPR31[17] ), .Y(
        OR4_29_Y));
    OR4 \OR4_R_DATA[16]  (.A(OR4_330_Y), .B(OR4_6_Y), .C(OR4_129_Y), 
        .D(OR4_173_Y), .Y(R_DATA_c[16]));
    OR4 OR4_280 (.A(OR4_629_Y), .B(OR4_407_Y), .C(OR4_446_Y), .D(
        OR4_579_Y), .Y(OR4_280_Y));
    OR4 OR4_587 (.A(\Z\R_DATA_TEMPR16[48] ), .B(\Z\R_DATA_TEMPR17[48] )
        , .C(\Z\R_DATA_TEMPR18[48] ), .D(\Z\R_DATA_TEMPR19[48] ), .Y(
        OR4_587_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%27%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C1 (
        .A_DOUT({\Z\R_DATA_TEMPR27[79] , \Z\R_DATA_TEMPR27[78] , 
        \Z\R_DATA_TEMPR27[77] , \Z\R_DATA_TEMPR27[76] , 
        \Z\R_DATA_TEMPR27[75] , \Z\R_DATA_TEMPR27[74] , 
        \Z\R_DATA_TEMPR27[73] , \Z\R_DATA_TEMPR27[72] , 
        \Z\R_DATA_TEMPR27[71] , \Z\R_DATA_TEMPR27[70] , 
        \Z\R_DATA_TEMPR27[69] , \Z\R_DATA_TEMPR27[68] , 
        \Z\R_DATA_TEMPR27[67] , \Z\R_DATA_TEMPR27[66] , 
        \Z\R_DATA_TEMPR27[65] , \Z\R_DATA_TEMPR27[64] , 
        \Z\R_DATA_TEMPR27[63] , \Z\R_DATA_TEMPR27[62] , 
        \Z\R_DATA_TEMPR27[61] , \Z\R_DATA_TEMPR27[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR27[59] , \Z\R_DATA_TEMPR27[58] , 
        \Z\R_DATA_TEMPR27[57] , \Z\R_DATA_TEMPR27[56] , 
        \Z\R_DATA_TEMPR27[55] , \Z\R_DATA_TEMPR27[54] , 
        \Z\R_DATA_TEMPR27[53] , \Z\R_DATA_TEMPR27[52] , 
        \Z\R_DATA_TEMPR27[51] , \Z\R_DATA_TEMPR27[50] , 
        \Z\R_DATA_TEMPR27[49] , \Z\R_DATA_TEMPR27[48] , 
        \Z\R_DATA_TEMPR27[47] , \Z\R_DATA_TEMPR27[46] , 
        \Z\R_DATA_TEMPR27[45] , \Z\R_DATA_TEMPR27[44] , 
        \Z\R_DATA_TEMPR27[43] , \Z\R_DATA_TEMPR27[42] , 
        \Z\R_DATA_TEMPR27[41] , \Z\R_DATA_TEMPR27[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[27][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[6] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[6] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_545 (.A(\Z\R_DATA_TEMPR8[47] ), .B(\Z\R_DATA_TEMPR9[47] ), 
        .C(\Z\R_DATA_TEMPR10[47] ), .D(\Z\R_DATA_TEMPR11[47] ), .Y(
        OR4_545_Y));
    OR4 OR4_233 (.A(OR4_390_Y), .B(OR2_20_Y), .C(
        \Z\R_DATA_TEMPR22[66] ), .D(\Z\R_DATA_TEMPR23[66] ), .Y(
        OR4_233_Y));
    OR4 \OR4_R_DATA[41]  (.A(OR4_378_Y), .B(OR4_341_Y), .C(OR4_352_Y), 
        .D(OR4_120_Y), .Y(R_DATA_c[41]));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%3%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0 (
        .A_DOUT({\Z\R_DATA_TEMPR3[39] , \Z\R_DATA_TEMPR3[38] , 
        \Z\R_DATA_TEMPR3[37] , \Z\R_DATA_TEMPR3[36] , 
        \Z\R_DATA_TEMPR3[35] , \Z\R_DATA_TEMPR3[34] , 
        \Z\R_DATA_TEMPR3[33] , \Z\R_DATA_TEMPR3[32] , 
        \Z\R_DATA_TEMPR3[31] , \Z\R_DATA_TEMPR3[30] , 
        \Z\R_DATA_TEMPR3[29] , \Z\R_DATA_TEMPR3[28] , 
        \Z\R_DATA_TEMPR3[27] , \Z\R_DATA_TEMPR3[26] , 
        \Z\R_DATA_TEMPR3[25] , \Z\R_DATA_TEMPR3[24] , 
        \Z\R_DATA_TEMPR3[23] , \Z\R_DATA_TEMPR3[22] , 
        \Z\R_DATA_TEMPR3[21] , \Z\R_DATA_TEMPR3[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR3[19] , \Z\R_DATA_TEMPR3[18] , 
        \Z\R_DATA_TEMPR3[17] , \Z\R_DATA_TEMPR3[16] , 
        \Z\R_DATA_TEMPR3[15] , \Z\R_DATA_TEMPR3[14] , 
        \Z\R_DATA_TEMPR3[13] , \Z\R_DATA_TEMPR3[12] , 
        \Z\R_DATA_TEMPR3[11] , \Z\R_DATA_TEMPR3[10] , 
        \Z\R_DATA_TEMPR3[9] , \Z\R_DATA_TEMPR3[8] , 
        \Z\R_DATA_TEMPR3[7] , \Z\R_DATA_TEMPR3[6] , 
        \Z\R_DATA_TEMPR3[5] , \Z\R_DATA_TEMPR3[4] , 
        \Z\R_DATA_TEMPR3[3] , \Z\R_DATA_TEMPR3[2] , 
        \Z\R_DATA_TEMPR3[1] , \Z\R_DATA_TEMPR3[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[3][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[0] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[0] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_562 (.A(OR4_506_Y), .B(OR4_351_Y), .C(OR4_513_Y), .D(
        OR4_109_Y), .Y(OR4_562_Y));
    OR4 OR4_689 (.A(OR4_467_Y), .B(OR4_313_Y), .C(OR4_212_Y), .D(
        OR4_244_Y), .Y(OR4_689_Y));
    OR4 OR4_643 (.A(\Z\R_DATA_TEMPR4[51] ), .B(\Z\R_DATA_TEMPR5[51] ), 
        .C(\Z\R_DATA_TEMPR6[51] ), .D(\Z\R_DATA_TEMPR7[51] ), .Y(
        OR4_643_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%12%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0 (
        .A_DOUT({\Z\R_DATA_TEMPR12[39] , \Z\R_DATA_TEMPR12[38] , 
        \Z\R_DATA_TEMPR12[37] , \Z\R_DATA_TEMPR12[36] , 
        \Z\R_DATA_TEMPR12[35] , \Z\R_DATA_TEMPR12[34] , 
        \Z\R_DATA_TEMPR12[33] , \Z\R_DATA_TEMPR12[32] , 
        \Z\R_DATA_TEMPR12[31] , \Z\R_DATA_TEMPR12[30] , 
        \Z\R_DATA_TEMPR12[29] , \Z\R_DATA_TEMPR12[28] , 
        \Z\R_DATA_TEMPR12[27] , \Z\R_DATA_TEMPR12[26] , 
        \Z\R_DATA_TEMPR12[25] , \Z\R_DATA_TEMPR12[24] , 
        \Z\R_DATA_TEMPR12[23] , \Z\R_DATA_TEMPR12[22] , 
        \Z\R_DATA_TEMPR12[21] , \Z\R_DATA_TEMPR12[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR12[19] , \Z\R_DATA_TEMPR12[18] , 
        \Z\R_DATA_TEMPR12[17] , \Z\R_DATA_TEMPR12[16] , 
        \Z\R_DATA_TEMPR12[15] , \Z\R_DATA_TEMPR12[14] , 
        \Z\R_DATA_TEMPR12[13] , \Z\R_DATA_TEMPR12[12] , 
        \Z\R_DATA_TEMPR12[11] , \Z\R_DATA_TEMPR12[10] , 
        \Z\R_DATA_TEMPR12[9] , \Z\R_DATA_TEMPR12[8] , 
        \Z\R_DATA_TEMPR12[7] , \Z\R_DATA_TEMPR12[6] , 
        \Z\R_DATA_TEMPR12[5] , \Z\R_DATA_TEMPR12[4] , 
        \Z\R_DATA_TEMPR12[3] , \Z\R_DATA_TEMPR12[2] , 
        \Z\R_DATA_TEMPR12[1] , \Z\R_DATA_TEMPR12[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[12][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[3] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[3] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_286 (.A(OR4_606_Y), .B(OR2_7_Y), .C(\Z\R_DATA_TEMPR22[69] )
        , .D(\Z\R_DATA_TEMPR23[69] ), .Y(OR4_286_Y));
    OR4 OR4_78 (.A(\Z\R_DATA_TEMPR0[4] ), .B(\Z\R_DATA_TEMPR1[4] ), .C(
        \Z\R_DATA_TEMPR2[4] ), .D(\Z\R_DATA_TEMPR3[4] ), .Y(OR4_78_Y));
    OR4 \OR4_R_DATA[8]  (.A(OR4_362_Y), .B(OR4_441_Y), .C(OR4_275_Y), 
        .D(OR4_542_Y), .Y(R_DATA_c[8]));
    OR4 \OR4_R_DATA[40]  (.A(OR4_256_Y), .B(OR4_403_Y), .C(OR4_10_Y), 
        .D(OR4_454_Y), .Y(R_DATA_c[40]));
    OR4 OR4_564 (.A(OR4_190_Y), .B(OR2_1_Y), .C(\Z\R_DATA_TEMPR22[78] )
        , .D(\Z\R_DATA_TEMPR23[78] ), .Y(OR4_564_Y));
    OR4 \OR4_R_DATA[61]  (.A(OR4_230_Y), .B(OR4_193_Y), .C(OR4_210_Y), 
        .D(OR4_697_Y), .Y(R_DATA_c[61]));
    OR4 OR4_154 (.A(OR4_223_Y), .B(OR4_614_Y), .C(OR4_167_Y), .D(
        OR4_512_Y), .Y(OR4_154_Y));
    OR4 OR4_684 (.A(\Z\R_DATA_TEMPR0[16] ), .B(\Z\R_DATA_TEMPR1[16] ), 
        .C(\Z\R_DATA_TEMPR2[16] ), .D(\Z\R_DATA_TEMPR3[16] ), .Y(
        OR4_684_Y));
    OR2 OR2_21 (.A(\Z\R_DATA_TEMPR20[3] ), .B(\Z\R_DATA_TEMPR21[3] ), 
        .Y(OR2_21_Y));
    OR4 OR4_638 (.A(\Z\R_DATA_TEMPR0[38] ), .B(\Z\R_DATA_TEMPR1[38] ), 
        .C(\Z\R_DATA_TEMPR2[38] ), .D(\Z\R_DATA_TEMPR3[38] ), .Y(
        OR4_638_Y));
    OR4 OR4_22 (.A(\Z\R_DATA_TEMPR8[41] ), .B(\Z\R_DATA_TEMPR9[41] ), 
        .C(\Z\R_DATA_TEMPR10[41] ), .D(\Z\R_DATA_TEMPR11[41] ), .Y(
        OR4_22_Y));
    OR2 OR2_73 (.A(\Z\R_DATA_TEMPR20[75] ), .B(\Z\R_DATA_TEMPR21[75] ), 
        .Y(OR2_73_Y));
    OR4 \OR4_R_DATA[46]  (.A(OR4_713_Y), .B(OR4_381_Y), .C(OR4_510_Y), 
        .D(OR4_548_Y), .Y(R_DATA_c[46]));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%29%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0 (
        .A_DOUT({\Z\R_DATA_TEMPR29[39] , \Z\R_DATA_TEMPR29[38] , 
        \Z\R_DATA_TEMPR29[37] , \Z\R_DATA_TEMPR29[36] , 
        \Z\R_DATA_TEMPR29[35] , \Z\R_DATA_TEMPR29[34] , 
        \Z\R_DATA_TEMPR29[33] , \Z\R_DATA_TEMPR29[32] , 
        \Z\R_DATA_TEMPR29[31] , \Z\R_DATA_TEMPR29[30] , 
        \Z\R_DATA_TEMPR29[29] , \Z\R_DATA_TEMPR29[28] , 
        \Z\R_DATA_TEMPR29[27] , \Z\R_DATA_TEMPR29[26] , 
        \Z\R_DATA_TEMPR29[25] , \Z\R_DATA_TEMPR29[24] , 
        \Z\R_DATA_TEMPR29[23] , \Z\R_DATA_TEMPR29[22] , 
        \Z\R_DATA_TEMPR29[21] , \Z\R_DATA_TEMPR29[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR29[19] , \Z\R_DATA_TEMPR29[18] , 
        \Z\R_DATA_TEMPR29[17] , \Z\R_DATA_TEMPR29[16] , 
        \Z\R_DATA_TEMPR29[15] , \Z\R_DATA_TEMPR29[14] , 
        \Z\R_DATA_TEMPR29[13] , \Z\R_DATA_TEMPR29[12] , 
        \Z\R_DATA_TEMPR29[11] , \Z\R_DATA_TEMPR29[10] , 
        \Z\R_DATA_TEMPR29[9] , \Z\R_DATA_TEMPR29[8] , 
        \Z\R_DATA_TEMPR29[7] , \Z\R_DATA_TEMPR29[6] , 
        \Z\R_DATA_TEMPR29[5] , \Z\R_DATA_TEMPR29[4] , 
        \Z\R_DATA_TEMPR29[3] , \Z\R_DATA_TEMPR29[2] , 
        \Z\R_DATA_TEMPR29[1] , \Z\R_DATA_TEMPR29[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[29][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[7] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[7] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_143 (.A(\Z\R_DATA_TEMPR12[8] ), .B(\Z\R_DATA_TEMPR13[8] ), 
        .C(\Z\R_DATA_TEMPR14[8] ), .D(\Z\R_DATA_TEMPR15[8] ), .Y(
        OR4_143_Y));
    OR4 OR4_632 (.A(\Z\R_DATA_TEMPR24[50] ), .B(\Z\R_DATA_TEMPR25[50] )
        , .C(\Z\R_DATA_TEMPR26[50] ), .D(\Z\R_DATA_TEMPR27[50] ), .Y(
        OR4_632_Y));
    OR4 OR4_213 (.A(\Z\R_DATA_TEMPR24[73] ), .B(\Z\R_DATA_TEMPR25[73] )
        , .C(\Z\R_DATA_TEMPR26[73] ), .D(\Z\R_DATA_TEMPR27[73] ), .Y(
        OR4_213_Y));
    OR4 OR4_201 (.A(\Z\R_DATA_TEMPR4[43] ), .B(\Z\R_DATA_TEMPR5[43] ), 
        .C(\Z\R_DATA_TEMPR6[43] ), .D(\Z\R_DATA_TEMPR7[43] ), .Y(
        OR4_201_Y));
    OR4 \OR4_R_DATA[74]  (.A(OR4_660_Y), .B(OR4_402_Y), .C(OR4_39_Y), 
        .D(OR4_348_Y), .Y(R_DATA_c[74]));
    OR4 OR4_361 (.A(\Z\R_DATA_TEMPR28[18] ), .B(\Z\R_DATA_TEMPR29[18] )
        , .C(\Z\R_DATA_TEMPR30[18] ), .D(\Z\R_DATA_TEMPR31[18] ), .Y(
        OR4_361_Y));
    OR4 \OR4_R_DATA[60]  (.A(OR4_81_Y), .B(OR4_263_Y), .C(OR4_578_Y), 
        .D(OR4_299_Y), .Y(R_DATA_c[60]));
    OR2 OR2_13 (.A(\Z\R_DATA_TEMPR20[5] ), .B(\Z\R_DATA_TEMPR21[5] ), 
        .Y(OR2_13_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%21%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0 (
        .A_DOUT({\Z\R_DATA_TEMPR21[39] , \Z\R_DATA_TEMPR21[38] , 
        \Z\R_DATA_TEMPR21[37] , \Z\R_DATA_TEMPR21[36] , 
        \Z\R_DATA_TEMPR21[35] , \Z\R_DATA_TEMPR21[34] , 
        \Z\R_DATA_TEMPR21[33] , \Z\R_DATA_TEMPR21[32] , 
        \Z\R_DATA_TEMPR21[31] , \Z\R_DATA_TEMPR21[30] , 
        \Z\R_DATA_TEMPR21[29] , \Z\R_DATA_TEMPR21[28] , 
        \Z\R_DATA_TEMPR21[27] , \Z\R_DATA_TEMPR21[26] , 
        \Z\R_DATA_TEMPR21[25] , \Z\R_DATA_TEMPR21[24] , 
        \Z\R_DATA_TEMPR21[23] , \Z\R_DATA_TEMPR21[22] , 
        \Z\R_DATA_TEMPR21[21] , \Z\R_DATA_TEMPR21[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR21[19] , \Z\R_DATA_TEMPR21[18] , 
        \Z\R_DATA_TEMPR21[17] , \Z\R_DATA_TEMPR21[16] , 
        \Z\R_DATA_TEMPR21[15] , \Z\R_DATA_TEMPR21[14] , 
        \Z\R_DATA_TEMPR21[13] , \Z\R_DATA_TEMPR21[12] , 
        \Z\R_DATA_TEMPR21[11] , \Z\R_DATA_TEMPR21[10] , 
        \Z\R_DATA_TEMPR21[9] , \Z\R_DATA_TEMPR21[8] , 
        \Z\R_DATA_TEMPR21[7] , \Z\R_DATA_TEMPR21[6] , 
        \Z\R_DATA_TEMPR21[5] , \Z\R_DATA_TEMPR21[4] , 
        \Z\R_DATA_TEMPR21[3] , \Z\R_DATA_TEMPR21[2] , 
        \Z\R_DATA_TEMPR21[1] , \Z\R_DATA_TEMPR21[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[21][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[5] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[5] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_6 (.A(OR4_182_Y), .B(OR2_67_Y), .C(\Z\R_DATA_TEMPR22[16] ), 
        .D(\Z\R_DATA_TEMPR23[16] ), .Y(OR4_6_Y));
    OR4 OR4_271 (.A(\Z\R_DATA_TEMPR4[45] ), .B(\Z\R_DATA_TEMPR5[45] ), 
        .C(\Z\R_DATA_TEMPR6[45] ), .D(\Z\R_DATA_TEMPR7[45] ), .Y(
        OR4_271_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%24%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C1 (
        .A_DOUT({\Z\R_DATA_TEMPR24[79] , \Z\R_DATA_TEMPR24[78] , 
        \Z\R_DATA_TEMPR24[77] , \Z\R_DATA_TEMPR24[76] , 
        \Z\R_DATA_TEMPR24[75] , \Z\R_DATA_TEMPR24[74] , 
        \Z\R_DATA_TEMPR24[73] , \Z\R_DATA_TEMPR24[72] , 
        \Z\R_DATA_TEMPR24[71] , \Z\R_DATA_TEMPR24[70] , 
        \Z\R_DATA_TEMPR24[69] , \Z\R_DATA_TEMPR24[68] , 
        \Z\R_DATA_TEMPR24[67] , \Z\R_DATA_TEMPR24[66] , 
        \Z\R_DATA_TEMPR24[65] , \Z\R_DATA_TEMPR24[64] , 
        \Z\R_DATA_TEMPR24[63] , \Z\R_DATA_TEMPR24[62] , 
        \Z\R_DATA_TEMPR24[61] , \Z\R_DATA_TEMPR24[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR24[59] , \Z\R_DATA_TEMPR24[58] , 
        \Z\R_DATA_TEMPR24[57] , \Z\R_DATA_TEMPR24[56] , 
        \Z\R_DATA_TEMPR24[55] , \Z\R_DATA_TEMPR24[54] , 
        \Z\R_DATA_TEMPR24[53] , \Z\R_DATA_TEMPR24[52] , 
        \Z\R_DATA_TEMPR24[51] , \Z\R_DATA_TEMPR24[50] , 
        \Z\R_DATA_TEMPR24[49] , \Z\R_DATA_TEMPR24[48] , 
        \Z\R_DATA_TEMPR24[47] , \Z\R_DATA_TEMPR24[46] , 
        \Z\R_DATA_TEMPR24[45] , \Z\R_DATA_TEMPR24[44] , 
        \Z\R_DATA_TEMPR24[43] , \Z\R_DATA_TEMPR24[42] , 
        \Z\R_DATA_TEMPR24[41] , \Z\R_DATA_TEMPR24[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[24][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[6] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[6] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_460 (.A(\Z\R_DATA_TEMPR12[63] ), .B(\Z\R_DATA_TEMPR13[63] )
        , .C(\Z\R_DATA_TEMPR14[63] ), .D(\Z\R_DATA_TEMPR15[63] ), .Y(
        OR4_460_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%28%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0 (
        .A_DOUT({\Z\R_DATA_TEMPR28[39] , \Z\R_DATA_TEMPR28[38] , 
        \Z\R_DATA_TEMPR28[37] , \Z\R_DATA_TEMPR28[36] , 
        \Z\R_DATA_TEMPR28[35] , \Z\R_DATA_TEMPR28[34] , 
        \Z\R_DATA_TEMPR28[33] , \Z\R_DATA_TEMPR28[32] , 
        \Z\R_DATA_TEMPR28[31] , \Z\R_DATA_TEMPR28[30] , 
        \Z\R_DATA_TEMPR28[29] , \Z\R_DATA_TEMPR28[28] , 
        \Z\R_DATA_TEMPR28[27] , \Z\R_DATA_TEMPR28[26] , 
        \Z\R_DATA_TEMPR28[25] , \Z\R_DATA_TEMPR28[24] , 
        \Z\R_DATA_TEMPR28[23] , \Z\R_DATA_TEMPR28[22] , 
        \Z\R_DATA_TEMPR28[21] , \Z\R_DATA_TEMPR28[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR28[19] , \Z\R_DATA_TEMPR28[18] , 
        \Z\R_DATA_TEMPR28[17] , \Z\R_DATA_TEMPR28[16] , 
        \Z\R_DATA_TEMPR28[15] , \Z\R_DATA_TEMPR28[14] , 
        \Z\R_DATA_TEMPR28[13] , \Z\R_DATA_TEMPR28[12] , 
        \Z\R_DATA_TEMPR28[11] , \Z\R_DATA_TEMPR28[10] , 
        \Z\R_DATA_TEMPR28[9] , \Z\R_DATA_TEMPR28[8] , 
        \Z\R_DATA_TEMPR28[7] , \Z\R_DATA_TEMPR28[6] , 
        \Z\R_DATA_TEMPR28[5] , \Z\R_DATA_TEMPR28[4] , 
        \Z\R_DATA_TEMPR28[3] , \Z\R_DATA_TEMPR28[2] , 
        \Z\R_DATA_TEMPR28[1] , \Z\R_DATA_TEMPR28[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[28][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[7] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[7] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[66]  (.A(OR4_558_Y), .B(OR4_233_Y), .C(OR4_350_Y), 
        .D(OR4_388_Y), .Y(R_DATA_c[66]));
    OR4 OR4_502 (.A(OR4_209_Y), .B(OR2_4_Y), .C(\Z\R_DATA_TEMPR22[12] )
        , .D(\Z\R_DATA_TEMPR23[12] ), .Y(OR4_502_Y));
    OR4 OR4_556 (.A(OR4_78_Y), .B(OR4_225_Y), .C(OR4_86_Y), .D(
        OR4_463_Y), .Y(OR4_556_Y));
    OR4 OR4_495 (.A(OR4_626_Y), .B(OR4_322_Y), .C(OR4_486_Y), .D(
        OR4_108_Y), .Y(OR4_495_Y));
    OR4 OR4_572 (.A(\Z\R_DATA_TEMPR0[14] ), .B(\Z\R_DATA_TEMPR1[14] ), 
        .C(\Z\R_DATA_TEMPR2[14] ), .D(\Z\R_DATA_TEMPR3[14] ), .Y(
        OR4_572_Y));
    OR2 OR2_54 (.A(\Z\R_DATA_TEMPR20[59] ), .B(\Z\R_DATA_TEMPR21[59] ), 
        .Y(OR2_54_Y));
    OR4 OR4_618 (.A(\Z\R_DATA_TEMPR24[62] ), .B(\Z\R_DATA_TEMPR25[62] )
        , .C(\Z\R_DATA_TEMPR26[62] ), .D(\Z\R_DATA_TEMPR27[62] ), .Y(
        OR4_618_Y));
    OR2 OR2_71 (.A(\Z\R_DATA_TEMPR20[27] ), .B(\Z\R_DATA_TEMPR21[27] ), 
        .Y(OR2_71_Y));
    OR4 \OR4_R_DATA[17]  (.A(OR4_154_Y), .B(OR4_501_Y), .C(OR4_682_Y), 
        .D(OR4_29_Y), .Y(R_DATA_c[17]));
    OR4 OR4_142 (.A(\Z\R_DATA_TEMPR24[31] ), .B(\Z\R_DATA_TEMPR25[31] )
        , .C(\Z\R_DATA_TEMPR26[31] ), .D(\Z\R_DATA_TEMPR27[31] ), .Y(
        OR4_142_Y));
    OR4 OR4_612 (.A(\Z\R_DATA_TEMPR4[15] ), .B(\Z\R_DATA_TEMPR5[15] ), 
        .C(\Z\R_DATA_TEMPR6[15] ), .D(\Z\R_DATA_TEMPR7[15] ), .Y(
        OR4_612_Y));
    OR4 OR4_504 (.A(OR4_121_Y), .B(OR4_644_Y), .C(OR4_676_Y), .D(
        OR4_73_Y), .Y(OR4_504_Y));
    OR4 OR4_574 (.A(\Z\R_DATA_TEMPR8[48] ), .B(\Z\R_DATA_TEMPR9[48] ), 
        .C(\Z\R_DATA_TEMPR10[48] ), .D(\Z\R_DATA_TEMPR11[48] ), .Y(
        OR4_574_Y));
    OR2 OR2_11 (.A(\Z\R_DATA_TEMPR20[50] ), .B(\Z\R_DATA_TEMPR21[50] ), 
        .Y(OR2_11_Y));
    OR4 OR4_494 (.A(\Z\R_DATA_TEMPR28[35] ), .B(\Z\R_DATA_TEMPR29[35] )
        , .C(\Z\R_DATA_TEMPR30[35] ), .D(\Z\R_DATA_TEMPR31[35] ), .Y(
        OR4_494_Y));
    OR4 OR4_558 (.A(OR4_188_Y), .B(OR4_687_Y), .C(OR4_1_Y), .D(
        OR4_124_Y), .Y(OR4_558_Y));
    OR4 OR4_55 (.A(\Z\R_DATA_TEMPR12[57] ), .B(\Z\R_DATA_TEMPR13[57] ), 
        .C(\Z\R_DATA_TEMPR14[57] ), .D(\Z\R_DATA_TEMPR15[57] ), .Y(
        OR4_55_Y));
    OR4 OR4_369 (.A(OR4_426_Y), .B(OR4_95_Y), .C(OR4_385_Y), .D(
        OR4_5_Y), .Y(OR4_369_Y));
    OR4 OR4_301 (.A(\Z\R_DATA_TEMPR24[20] ), .B(\Z\R_DATA_TEMPR25[20] )
        , .C(\Z\R_DATA_TEMPR26[20] ), .D(\Z\R_DATA_TEMPR27[20] ), .Y(
        OR4_301_Y));
    OR4 OR4_396 (.A(\Z\R_DATA_TEMPR12[38] ), .B(\Z\R_DATA_TEMPR13[38] )
        , .C(\Z\R_DATA_TEMPR14[38] ), .D(\Z\R_DATA_TEMPR15[38] ), .Y(
        OR4_396_Y));
    OR4 OR4_249 (.A(OR4_12_Y), .B(OR4_588_Y), .C(OR4_465_Y), .D(
        OR4_500_Y), .Y(OR4_249_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%1%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0 (
        .A_DOUT({\Z\R_DATA_TEMPR1[39] , \Z\R_DATA_TEMPR1[38] , 
        \Z\R_DATA_TEMPR1[37] , \Z\R_DATA_TEMPR1[36] , 
        \Z\R_DATA_TEMPR1[35] , \Z\R_DATA_TEMPR1[34] , 
        \Z\R_DATA_TEMPR1[33] , \Z\R_DATA_TEMPR1[32] , 
        \Z\R_DATA_TEMPR1[31] , \Z\R_DATA_TEMPR1[30] , 
        \Z\R_DATA_TEMPR1[29] , \Z\R_DATA_TEMPR1[28] , 
        \Z\R_DATA_TEMPR1[27] , \Z\R_DATA_TEMPR1[26] , 
        \Z\R_DATA_TEMPR1[25] , \Z\R_DATA_TEMPR1[24] , 
        \Z\R_DATA_TEMPR1[23] , \Z\R_DATA_TEMPR1[22] , 
        \Z\R_DATA_TEMPR1[21] , \Z\R_DATA_TEMPR1[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR1[19] , \Z\R_DATA_TEMPR1[18] , 
        \Z\R_DATA_TEMPR1[17] , \Z\R_DATA_TEMPR1[16] , 
        \Z\R_DATA_TEMPR1[15] , \Z\R_DATA_TEMPR1[14] , 
        \Z\R_DATA_TEMPR1[13] , \Z\R_DATA_TEMPR1[12] , 
        \Z\R_DATA_TEMPR1[11] , \Z\R_DATA_TEMPR1[10] , 
        \Z\R_DATA_TEMPR1[9] , \Z\R_DATA_TEMPR1[8] , 
        \Z\R_DATA_TEMPR1[7] , \Z\R_DATA_TEMPR1[6] , 
        \Z\R_DATA_TEMPR1[5] , \Z\R_DATA_TEMPR1[4] , 
        \Z\R_DATA_TEMPR1[3] , \Z\R_DATA_TEMPR1[2] , 
        \Z\R_DATA_TEMPR1[1] , \Z\R_DATA_TEMPR1[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[1][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[0] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[0] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_425 (.A(\Z\R_DATA_TEMPR24[38] ), .B(\Z\R_DATA_TEMPR25[38] )
        , .C(\Z\R_DATA_TEMPR26[38] ), .D(\Z\R_DATA_TEMPR27[38] ), .Y(
        OR4_425_Y));
    OR4 OR4_371 (.A(\Z\R_DATA_TEMPR28[3] ), .B(\Z\R_DATA_TEMPR29[3] ), 
        .C(\Z\R_DATA_TEMPR30[3] ), .D(\Z\R_DATA_TEMPR31[3] ), .Y(
        OR4_371_Y));
    OR4 OR4_400 (.A(\Z\R_DATA_TEMPR28[47] ), .B(\Z\R_DATA_TEMPR29[47] )
        , .C(\Z\R_DATA_TEMPR30[47] ), .D(\Z\R_DATA_TEMPR31[47] ), .Y(
        OR4_400_Y));
    OR4 \OR4_R_DATA[38]  (.A(OR4_125_Y), .B(OR4_38_Y), .C(OR4_425_Y), 
        .D(OR4_531_Y), .Y(R_DATA_c[38]));
    OR4 OR4_636 (.A(OR4_204_Y), .B(OR4_612_Y), .C(OR4_646_Y), .D(
        OR4_284_Y), .Y(OR4_636_Y));
    OR4 OR4_456 (.A(\Z\R_DATA_TEMPR0[55] ), .B(\Z\R_DATA_TEMPR1[55] ), 
        .C(\Z\R_DATA_TEMPR2[55] ), .D(\Z\R_DATA_TEMPR3[55] ), .Y(
        OR4_456_Y));
    OR4 OR4_470 (.A(\Z\R_DATA_TEMPR28[53] ), .B(\Z\R_DATA_TEMPR29[53] )
        , .C(\Z\R_DATA_TEMPR30[53] ), .D(\Z\R_DATA_TEMPR31[53] ), .Y(
        OR4_470_Y));
    OR4 \OR4_R_DATA[47]  (.A(OR4_530_Y), .B(OR4_153_Y), .C(OR4_329_Y), 
        .D(OR4_400_Y), .Y(R_DATA_c[47]));
    OR4 OR4_352 (.A(\Z\R_DATA_TEMPR24[41] ), .B(\Z\R_DATA_TEMPR25[41] )
        , .C(\Z\R_DATA_TEMPR26[41] ), .D(\Z\R_DATA_TEMPR27[41] ), .Y(
        OR4_352_Y));
    OR4 OR4_15 (.A(\Z\R_DATA_TEMPR0[69] ), .B(\Z\R_DATA_TEMPR1[69] ), 
        .C(\Z\R_DATA_TEMPR2[69] ), .D(\Z\R_DATA_TEMPR3[69] ), .Y(
        OR4_15_Y));
    GND GND_Z (.Y(GND));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKX2[3]  (.A(CFG2_0_Y), .B(
        W_ADDR_c[13]), .C(W_EN_c), .Y(\Z\BLKX2[3] ));
    OR4 OR4_424 (.A(\Z\R_DATA_TEMPR16[68] ), .B(\Z\R_DATA_TEMPR17[68] )
        , .C(\Z\R_DATA_TEMPR18[68] ), .D(\Z\R_DATA_TEMPR19[68] ), .Y(
        OR4_424_Y));
    OR4 OR4_281 (.A(\Z\R_DATA_TEMPR16[44] ), .B(\Z\R_DATA_TEMPR17[44] )
        , .C(\Z\R_DATA_TEMPR18[44] ), .D(\Z\R_DATA_TEMPR19[44] ), .Y(
        OR4_281_Y));
    OR4 \OR4_R_DATA[67]  (.A(OR4_369_Y), .B(OR4_715_Y), .C(OR4_186_Y), 
        .D(OR4_257_Y), .Y(R_DATA_c[67]));
    OR4 OR4_326 (.A(\Z\R_DATA_TEMPR28[78] ), .B(\Z\R_DATA_TEMPR29[78] )
        , .C(\Z\R_DATA_TEMPR30[78] ), .D(\Z\R_DATA_TEMPR31[78] ), .Y(
        OR4_326_Y));
    OR4 OR4_194 (.A(\Z\R_DATA_TEMPR24[45] ), .B(\Z\R_DATA_TEMPR25[45] )
        , .C(\Z\R_DATA_TEMPR26[45] ), .D(\Z\R_DATA_TEMPR27[45] ), .Y(
        OR4_194_Y));
    OR4 OR4_93 (.A(\Z\R_DATA_TEMPR12[64] ), .B(\Z\R_DATA_TEMPR13[64] ), 
        .C(\Z\R_DATA_TEMPR14[64] ), .D(\Z\R_DATA_TEMPR15[64] ), .Y(
        OR4_93_Y));
    OR4 OR4_563 (.A(\Z\R_DATA_TEMPR16[37] ), .B(\Z\R_DATA_TEMPR17[37] )
        , .C(\Z\R_DATA_TEMPR18[37] ), .D(\Z\R_DATA_TEMPR19[37] ), .Y(
        OR4_563_Y));
    OR4 OR4_616 (.A(\Z\R_DATA_TEMPR16[67] ), .B(\Z\R_DATA_TEMPR17[67] )
        , .C(\Z\R_DATA_TEMPR18[67] ), .D(\Z\R_DATA_TEMPR19[67] ), .Y(
        OR4_616_Y));
    OR4 OR4_309 (.A(OR4_659_Y), .B(OR4_438_Y), .C(OR4_487_Y), .D(
        OR4_613_Y), .Y(OR4_309_Y));
    OR4 OR4_582 (.A(\Z\R_DATA_TEMPR8[25] ), .B(\Z\R_DATA_TEMPR9[25] ), 
        .C(\Z\R_DATA_TEMPR10[25] ), .D(\Z\R_DATA_TEMPR11[25] ), .Y(
        OR4_582_Y));
    OR4 OR4_24 (.A(\Z\R_DATA_TEMPR24[19] ), .B(\Z\R_DATA_TEMPR25[19] ), 
        .C(\Z\R_DATA_TEMPR26[19] ), .D(\Z\R_DATA_TEMPR27[19] ), .Y(
        OR4_24_Y));
    OR4 OR4_8 (.A(\Z\R_DATA_TEMPR4[42] ), .B(\Z\R_DATA_TEMPR5[42] ), 
        .C(\Z\R_DATA_TEMPR6[42] ), .D(\Z\R_DATA_TEMPR7[42] ), .Y(
        OR4_8_Y));
    OR4 OR4_379 (.A(\Z\R_DATA_TEMPR0[37] ), .B(\Z\R_DATA_TEMPR1[37] ), 
        .C(\Z\R_DATA_TEMPR2[37] ), .D(\Z\R_DATA_TEMPR3[37] ), .Y(
        OR4_379_Y));
    OR4 OR4_250 (.A(OR4_442_Y), .B(OR2_31_Y), .C(
        \Z\R_DATA_TEMPR22[51] ), .D(\Z\R_DATA_TEMPR23[51] ), .Y(
        OR4_250_Y));
    OR4 OR4_557 (.A(\Z\R_DATA_TEMPR12[55] ), .B(\Z\R_DATA_TEMPR13[55] )
        , .C(\Z\R_DATA_TEMPR14[55] ), .D(\Z\R_DATA_TEMPR15[55] ), .Y(
        OR4_557_Y));
    OR4 OR4_334 (.A(\Z\R_DATA_TEMPR0[46] ), .B(\Z\R_DATA_TEMPR1[46] ), 
        .C(\Z\R_DATA_TEMPR2[46] ), .D(\Z\R_DATA_TEMPR3[46] ), .Y(
        OR4_334_Y));
    OR2 OR2_4 (.A(\Z\R_DATA_TEMPR20[12] ), .B(\Z\R_DATA_TEMPR21[12] ), 
        .Y(OR2_4_Y));
    OR4 \OR4_R_DATA[71]  (.A(OR4_700_Y), .B(OR4_664_Y), .C(OR4_674_Y), 
        .D(OR4_447_Y), .Y(R_DATA_c[71]));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%18%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C1 (
        .A_DOUT({\Z\R_DATA_TEMPR18[79] , \Z\R_DATA_TEMPR18[78] , 
        \Z\R_DATA_TEMPR18[77] , \Z\R_DATA_TEMPR18[76] , 
        \Z\R_DATA_TEMPR18[75] , \Z\R_DATA_TEMPR18[74] , 
        \Z\R_DATA_TEMPR18[73] , \Z\R_DATA_TEMPR18[72] , 
        \Z\R_DATA_TEMPR18[71] , \Z\R_DATA_TEMPR18[70] , 
        \Z\R_DATA_TEMPR18[69] , \Z\R_DATA_TEMPR18[68] , 
        \Z\R_DATA_TEMPR18[67] , \Z\R_DATA_TEMPR18[66] , 
        \Z\R_DATA_TEMPR18[65] , \Z\R_DATA_TEMPR18[64] , 
        \Z\R_DATA_TEMPR18[63] , \Z\R_DATA_TEMPR18[62] , 
        \Z\R_DATA_TEMPR18[61] , \Z\R_DATA_TEMPR18[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR18[59] , \Z\R_DATA_TEMPR18[58] , 
        \Z\R_DATA_TEMPR18[57] , \Z\R_DATA_TEMPR18[56] , 
        \Z\R_DATA_TEMPR18[55] , \Z\R_DATA_TEMPR18[54] , 
        \Z\R_DATA_TEMPR18[53] , \Z\R_DATA_TEMPR18[52] , 
        \Z\R_DATA_TEMPR18[51] , \Z\R_DATA_TEMPR18[50] , 
        \Z\R_DATA_TEMPR18[49] , \Z\R_DATA_TEMPR18[48] , 
        \Z\R_DATA_TEMPR18[47] , \Z\R_DATA_TEMPR18[46] , 
        \Z\R_DATA_TEMPR18[45] , \Z\R_DATA_TEMPR18[44] , 
        \Z\R_DATA_TEMPR18[43] , \Z\R_DATA_TEMPR18[42] , 
        \Z\R_DATA_TEMPR18[41] , \Z\R_DATA_TEMPR18[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[18][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[4] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[4] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_131 (.A(OR4_72_Y), .B(OR4_651_Y), .C(OR4_79_Y), .D(
        OR4_414_Y), .Y(OR4_131_Y));
    OR4 OR4_584 (.A(\Z\R_DATA_TEMPR4[77] ), .B(\Z\R_DATA_TEMPR5[77] ), 
        .C(\Z\R_DATA_TEMPR6[77] ), .D(\Z\R_DATA_TEMPR7[77] ), .Y(
        OR4_584_Y));
    OR4 OR4_659 (.A(\Z\R_DATA_TEMPR0[76] ), .B(\Z\R_DATA_TEMPR1[76] ), 
        .C(\Z\R_DATA_TEMPR2[76] ), .D(\Z\R_DATA_TEMPR3[76] ), .Y(
        OR4_659_Y));
    OR4 OR4_596 (.A(\Z\R_DATA_TEMPR0[22] ), .B(\Z\R_DATA_TEMPR1[22] ), 
        .C(\Z\R_DATA_TEMPR2[22] ), .D(\Z\R_DATA_TEMPR3[22] ), .Y(
        OR4_596_Y));
    OR4 \OR4_R_DATA[39]  (.A(OR4_393_Y), .B(OR4_252_Y), .C(OR4_202_Y), 
        .D(OR4_58_Y), .Y(R_DATA_c[39]));
    OR4 OR4_256 (.A(OR4_199_Y), .B(OR4_35_Y), .C(OR4_207_Y), .D(
        OR4_523_Y), .Y(OR4_256_Y));
    OR2 OR2_0 (.A(\Z\R_DATA_TEMPR20[74] ), .B(\Z\R_DATA_TEMPR21[74] ), 
        .Y(OR2_0_Y));
    OR4 OR4_75 (.A(\Z\R_DATA_TEMPR4[53] ), .B(\Z\R_DATA_TEMPR5[53] ), 
        .C(\Z\R_DATA_TEMPR6[53] ), .D(\Z\R_DATA_TEMPR7[53] ), .Y(
        OR4_75_Y));
    OR2 OR2_6 (.A(\Z\R_DATA_TEMPR20[33] ), .B(\Z\R_DATA_TEMPR21[33] ), 
        .Y(OR2_6_Y));
    OR4 \OR4_R_DATA[70]  (.A(OR4_562_Y), .B(OR4_3_Y), .C(OR4_323_Y), 
        .D(OR4_54_Y), .Y(R_DATA_c[70]));
    OR4 OR4_431 (.A(\Z\R_DATA_TEMPR28[56] ), .B(\Z\R_DATA_TEMPR29[56] )
        , .C(\Z\R_DATA_TEMPR30[56] ), .D(\Z\R_DATA_TEMPR31[56] ), .Y(
        OR4_431_Y));
    OR4 OR4_91 (.A(\Z\R_DATA_TEMPR0[32] ), .B(\Z\R_DATA_TEMPR1[32] ), 
        .C(\Z\R_DATA_TEMPR2[32] ), .D(\Z\R_DATA_TEMPR3[32] ), .Y(
        OR4_91_Y));
    OR4 OR4_124 (.A(\Z\R_DATA_TEMPR12[66] ), .B(\Z\R_DATA_TEMPR13[66] )
        , .C(\Z\R_DATA_TEMPR14[66] ), .D(\Z\R_DATA_TEMPR15[66] ), .Y(
        OR4_124_Y));
    OR4 OR4_438 (.A(\Z\R_DATA_TEMPR4[76] ), .B(\Z\R_DATA_TEMPR5[76] ), 
        .C(\Z\R_DATA_TEMPR6[76] ), .D(\Z\R_DATA_TEMPR7[76] ), .Y(
        OR4_438_Y));
    OR4 OR4_709 (.A(\Z\R_DATA_TEMPR4[33] ), .B(\Z\R_DATA_TEMPR5[33] ), 
        .C(\Z\R_DATA_TEMPR6[33] ), .D(\Z\R_DATA_TEMPR7[33] ), .Y(
        OR4_709_Y));
    OR4 OR4_381 (.A(OR4_553_Y), .B(OR2_59_Y), .C(
        \Z\R_DATA_TEMPR22[46] ), .D(\Z\R_DATA_TEMPR23[46] ), .Y(
        OR4_381_Y));
    OR2 OR2_3 (.A(\Z\R_DATA_TEMPR20[71] ), .B(\Z\R_DATA_TEMPR21[71] ), 
        .Y(OR2_3_Y));
    OR4 OR4_654 (.A(\Z\R_DATA_TEMPR0[73] ), .B(\Z\R_DATA_TEMPR1[73] ), 
        .C(\Z\R_DATA_TEMPR2[73] ), .D(\Z\R_DATA_TEMPR3[73] ), .Y(
        OR4_654_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[5]  (.A(CFG2_2_Y), .B(
        W_ADDR_c[13]), .C(W_EN_c), .Y(\Z\BLKX2[5] ));
    OR4 \OR4_R_DATA[76]  (.A(OR4_309_Y), .B(OR4_705_Y), .C(OR4_97_Y), 
        .D(OR4_141_Y), .Y(R_DATA_c[76]));
    OR4 OR4_480 (.A(\Z\R_DATA_TEMPR24[1] ), .B(\Z\R_DATA_TEMPR25[1] ), 
        .C(\Z\R_DATA_TEMPR26[1] ), .D(\Z\R_DATA_TEMPR27[1] ), .Y(
        OR4_480_Y));
    OR4 OR4_503 (.A(\Z\R_DATA_TEMPR12[65] ), .B(\Z\R_DATA_TEMPR13[65] )
        , .C(\Z\R_DATA_TEMPR14[65] ), .D(\Z\R_DATA_TEMPR15[65] ), .Y(
        OR4_503_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[7]  (.A(CFG2_0_Y), .B(
        W_ADDR_c[13]), .C(W_EN_c), .Y(\Z\BLKX2[7] ));
    OR4 OR4_314 (.A(\Z\R_DATA_TEMPR24[3] ), .B(\Z\R_DATA_TEMPR25[3] ), 
        .C(\Z\R_DATA_TEMPR26[3] ), .D(\Z\R_DATA_TEMPR27[3] ), .Y(
        OR4_314_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%20%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0 (
        .A_DOUT({\Z\R_DATA_TEMPR20[39] , \Z\R_DATA_TEMPR20[38] , 
        \Z\R_DATA_TEMPR20[37] , \Z\R_DATA_TEMPR20[36] , 
        \Z\R_DATA_TEMPR20[35] , \Z\R_DATA_TEMPR20[34] , 
        \Z\R_DATA_TEMPR20[33] , \Z\R_DATA_TEMPR20[32] , 
        \Z\R_DATA_TEMPR20[31] , \Z\R_DATA_TEMPR20[30] , 
        \Z\R_DATA_TEMPR20[29] , \Z\R_DATA_TEMPR20[28] , 
        \Z\R_DATA_TEMPR20[27] , \Z\R_DATA_TEMPR20[26] , 
        \Z\R_DATA_TEMPR20[25] , \Z\R_DATA_TEMPR20[24] , 
        \Z\R_DATA_TEMPR20[23] , \Z\R_DATA_TEMPR20[22] , 
        \Z\R_DATA_TEMPR20[21] , \Z\R_DATA_TEMPR20[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR20[19] , \Z\R_DATA_TEMPR20[18] , 
        \Z\R_DATA_TEMPR20[17] , \Z\R_DATA_TEMPR20[16] , 
        \Z\R_DATA_TEMPR20[15] , \Z\R_DATA_TEMPR20[14] , 
        \Z\R_DATA_TEMPR20[13] , \Z\R_DATA_TEMPR20[12] , 
        \Z\R_DATA_TEMPR20[11] , \Z\R_DATA_TEMPR20[10] , 
        \Z\R_DATA_TEMPR20[9] , \Z\R_DATA_TEMPR20[8] , 
        \Z\R_DATA_TEMPR20[7] , \Z\R_DATA_TEMPR20[6] , 
        \Z\R_DATA_TEMPR20[5] , \Z\R_DATA_TEMPR20[4] , 
        \Z\R_DATA_TEMPR20[3] , \Z\R_DATA_TEMPR20[2] , 
        \Z\R_DATA_TEMPR20[1] , \Z\R_DATA_TEMPR20[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[20][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[5] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[5] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_43 (.A(OR4_668_Y), .B(OR2_45_Y), .C(\Z\R_DATA_TEMPR22[57] )
        , .D(\Z\R_DATA_TEMPR23[57] ), .Y(OR4_43_Y));
    OR4 OR4_573 (.A(\Z\R_DATA_TEMPR0[0] ), .B(\Z\R_DATA_TEMPR1[0] ), 
        .C(\Z\R_DATA_TEMPR2[0] ), .D(\Z\R_DATA_TEMPR3[0] ), .Y(
        OR4_573_Y));
    OR4 OR4_539 (.A(\Z\R_DATA_TEMPR0[10] ), .B(\Z\R_DATA_TEMPR1[10] ), 
        .C(\Z\R_DATA_TEMPR2[10] ), .D(\Z\R_DATA_TEMPR3[10] ), .Y(
        OR4_539_Y));
    OR4 OR4_111 (.A(\Z\R_DATA_TEMPR0[48] ), .B(\Z\R_DATA_TEMPR1[48] ), 
        .C(\Z\R_DATA_TEMPR2[48] ), .D(\Z\R_DATA_TEMPR3[48] ), .Y(
        OR4_111_Y));
    OR2 OR2_26 (.A(\Z\R_DATA_TEMPR20[54] ), .B(\Z\R_DATA_TEMPR21[54] ), 
        .Y(OR2_26_Y));
    INV \INVBLKX0[0]  (.A(W_ADDR_c[9]), .Y(\Z\BLKX0[0] ));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%16%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C1 (
        .A_DOUT({\Z\R_DATA_TEMPR16[79] , \Z\R_DATA_TEMPR16[78] , 
        \Z\R_DATA_TEMPR16[77] , \Z\R_DATA_TEMPR16[76] , 
        \Z\R_DATA_TEMPR16[75] , \Z\R_DATA_TEMPR16[74] , 
        \Z\R_DATA_TEMPR16[73] , \Z\R_DATA_TEMPR16[72] , 
        \Z\R_DATA_TEMPR16[71] , \Z\R_DATA_TEMPR16[70] , 
        \Z\R_DATA_TEMPR16[69] , \Z\R_DATA_TEMPR16[68] , 
        \Z\R_DATA_TEMPR16[67] , \Z\R_DATA_TEMPR16[66] , 
        \Z\R_DATA_TEMPR16[65] , \Z\R_DATA_TEMPR16[64] , 
        \Z\R_DATA_TEMPR16[63] , \Z\R_DATA_TEMPR16[62] , 
        \Z\R_DATA_TEMPR16[61] , \Z\R_DATA_TEMPR16[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR16[59] , \Z\R_DATA_TEMPR16[58] , 
        \Z\R_DATA_TEMPR16[57] , \Z\R_DATA_TEMPR16[56] , 
        \Z\R_DATA_TEMPR16[55] , \Z\R_DATA_TEMPR16[54] , 
        \Z\R_DATA_TEMPR16[53] , \Z\R_DATA_TEMPR16[52] , 
        \Z\R_DATA_TEMPR16[51] , \Z\R_DATA_TEMPR16[50] , 
        \Z\R_DATA_TEMPR16[49] , \Z\R_DATA_TEMPR16[48] , 
        \Z\R_DATA_TEMPR16[47] , \Z\R_DATA_TEMPR16[46] , 
        \Z\R_DATA_TEMPR16[45] , \Z\R_DATA_TEMPR16[44] , 
        \Z\R_DATA_TEMPR16[43] , \Z\R_DATA_TEMPR16[42] , 
        \Z\R_DATA_TEMPR16[41] , \Z\R_DATA_TEMPR16[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[16][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[4] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[4] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_598 (.A(\Z\R_DATA_TEMPR28[64] ), .B(\Z\R_DATA_TEMPR29[64] )
        , .C(\Z\R_DATA_TEMPR30[64] ), .D(\Z\R_DATA_TEMPR31[64] ), .Y(
        OR4_598_Y));
    OR4 OR4_59 (.A(\Z\R_DATA_TEMPR0[64] ), .B(\Z\R_DATA_TEMPR1[64] ), 
        .C(\Z\R_DATA_TEMPR2[64] ), .D(\Z\R_DATA_TEMPR3[64] ), .Y(
        OR4_59_Y));
    OR4 OR4_530 (.A(OR4_591_Y), .B(OR4_273_Y), .C(OR4_545_Y), .D(
        OR4_162_Y), .Y(OR4_530_Y));
    OR4 OR4_263 (.A(OR4_355_Y), .B(OR2_50_Y), .C(
        \Z\R_DATA_TEMPR22[60] ), .D(\Z\R_DATA_TEMPR23[60] ), .Y(
        OR4_263_Y));
    OR4 OR4_526 (.A(OR4_656_Y), .B(OR4_356_Y), .C(OR4_508_Y), .D(
        OR4_144_Y), .Y(OR4_526_Y));
    OR4 OR4_445 (.A(\Z\R_DATA_TEMPR8[22] ), .B(\Z\R_DATA_TEMPR9[22] ), 
        .C(\Z\R_DATA_TEMPR10[22] ), .D(\Z\R_DATA_TEMPR11[22] ), .Y(
        OR4_445_Y));
    OR4 OR4_411 (.A(\Z\R_DATA_TEMPR12[52] ), .B(\Z\R_DATA_TEMPR13[52] )
        , .C(\Z\R_DATA_TEMPR14[52] ), .D(\Z\R_DATA_TEMPR15[52] ), .Y(
        OR4_411_Y));
    OR4 OR4_496 (.A(\Z\R_DATA_TEMPR16[43] ), .B(\Z\R_DATA_TEMPR17[43] )
        , .C(\Z\R_DATA_TEMPR18[43] ), .D(\Z\R_DATA_TEMPR19[43] ), .Y(
        OR4_496_Y));
    OR4 OR4_418 (.A(OR4_130_Y), .B(OR2_30_Y), .C(
        \Z\R_DATA_TEMPR22[35] ), .D(\Z\R_DATA_TEMPR23[35] ), .Y(
        OR4_418_Y));
    OR4 \OR4_R_DATA[0]  (.A(OR4_599_Y), .B(OR4_680_Y), .C(OR4_452_Y), 
        .D(OR4_592_Y), .Y(R_DATA_c[0]));
    OR4 OR4_389 (.A(\Z\R_DATA_TEMPR16[53] ), .B(\Z\R_DATA_TEMPR17[53] )
        , .C(\Z\R_DATA_TEMPR18[53] ), .D(\Z\R_DATA_TEMPR19[53] ), .Y(
        OR4_389_Y));
    OR4 OR4_392 (.A(OR4_474_Y), .B(OR4_231_Y), .C(OR4_478_Y), .D(
        OR4_215_Y), .Y(OR4_392_Y));
    OR4 OR4_19 (.A(OR4_147_Y), .B(OR4_576_Y), .C(OR4_0_Y), .D(
        OR4_363_Y), .Y(OR4_19_Y));
    OR4 OR4_41 (.A(\Z\R_DATA_TEMPR16[49] ), .B(\Z\R_DATA_TEMPR17[49] ), 
        .C(\Z\R_DATA_TEMPR18[49] ), .D(\Z\R_DATA_TEMPR19[49] ), .Y(
        OR4_41_Y));
    OR4 OR4_333 (.A(\Z\R_DATA_TEMPR16[63] ), .B(\Z\R_DATA_TEMPR17[63] )
        , .C(\Z\R_DATA_TEMPR18[63] ), .D(\Z\R_DATA_TEMPR19[63] ), .Y(
        OR4_333_Y));
    OR4 OR4_519 (.A(\Z\R_DATA_TEMPR8[39] ), .B(\Z\R_DATA_TEMPR9[39] ), 
        .C(\Z\R_DATA_TEMPR10[39] ), .D(\Z\R_DATA_TEMPR11[39] ), .Y(
        OR4_519_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%17%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C1 (
        .A_DOUT({\Z\R_DATA_TEMPR17[79] , \Z\R_DATA_TEMPR17[78] , 
        \Z\R_DATA_TEMPR17[77] , \Z\R_DATA_TEMPR17[76] , 
        \Z\R_DATA_TEMPR17[75] , \Z\R_DATA_TEMPR17[74] , 
        \Z\R_DATA_TEMPR17[73] , \Z\R_DATA_TEMPR17[72] , 
        \Z\R_DATA_TEMPR17[71] , \Z\R_DATA_TEMPR17[70] , 
        \Z\R_DATA_TEMPR17[69] , \Z\R_DATA_TEMPR17[68] , 
        \Z\R_DATA_TEMPR17[67] , \Z\R_DATA_TEMPR17[66] , 
        \Z\R_DATA_TEMPR17[65] , \Z\R_DATA_TEMPR17[64] , 
        \Z\R_DATA_TEMPR17[63] , \Z\R_DATA_TEMPR17[62] , 
        \Z\R_DATA_TEMPR17[61] , \Z\R_DATA_TEMPR17[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR17[59] , \Z\R_DATA_TEMPR17[58] , 
        \Z\R_DATA_TEMPR17[57] , \Z\R_DATA_TEMPR17[56] , 
        \Z\R_DATA_TEMPR17[55] , \Z\R_DATA_TEMPR17[54] , 
        \Z\R_DATA_TEMPR17[53] , \Z\R_DATA_TEMPR17[52] , 
        \Z\R_DATA_TEMPR17[51] , \Z\R_DATA_TEMPR17[50] , 
        \Z\R_DATA_TEMPR17[49] , \Z\R_DATA_TEMPR17[48] , 
        \Z\R_DATA_TEMPR17[47] , \Z\R_DATA_TEMPR17[46] , 
        \Z\R_DATA_TEMPR17[45] , \Z\R_DATA_TEMPR17[44] , 
        \Z\R_DATA_TEMPR17[43] , \Z\R_DATA_TEMPR17[42] , 
        \Z\R_DATA_TEMPR17[41] , \Z\R_DATA_TEMPR17[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[17][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[4] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[4] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_668 (.A(\Z\R_DATA_TEMPR16[57] ), .B(\Z\R_DATA_TEMPR17[57] )
        , .C(\Z\R_DATA_TEMPR18[57] ), .D(\Z\R_DATA_TEMPR19[57] ), .Y(
        OR4_668_Y));
    OR4 OR4_510 (.A(\Z\R_DATA_TEMPR24[46] ), .B(\Z\R_DATA_TEMPR25[46] )
        , .C(\Z\R_DATA_TEMPR26[46] ), .D(\Z\R_DATA_TEMPR27[46] ), .Y(
        OR4_510_Y));
    OR4 OR4_444 (.A(\Z\R_DATA_TEMPR12[68] ), .B(\Z\R_DATA_TEMPR13[68] )
        , .C(\Z\R_DATA_TEMPR14[68] ), .D(\Z\R_DATA_TEMPR15[68] ), .Y(
        OR4_444_Y));
    OR4 OR4_432 (.A(\Z\R_DATA_TEMPR0[78] ), .B(\Z\R_DATA_TEMPR1[78] ), 
        .C(\Z\R_DATA_TEMPR2[78] ), .D(\Z\R_DATA_TEMPR3[78] ), .Y(
        OR4_432_Y));
    OR4 OR4_528 (.A(\Z\R_DATA_TEMPR8[13] ), .B(\Z\R_DATA_TEMPR9[13] ), 
        .C(\Z\R_DATA_TEMPR10[13] ), .D(\Z\R_DATA_TEMPR11[13] ), .Y(
        OR4_528_Y));
    OR4 OR4_52 (.A(\Z\R_DATA_TEMPR8[56] ), .B(\Z\R_DATA_TEMPR9[56] ), 
        .C(\Z\R_DATA_TEMPR10[56] ), .D(\Z\R_DATA_TEMPR11[56] ), .Y(
        OR4_52_Y));
    OR2 OR2_76 (.A(\Z\R_DATA_TEMPR20[13] ), .B(\Z\R_DATA_TEMPR21[13] ), 
        .Y(OR2_76_Y));
    OR4 OR4_662 (.A(OR4_432_Y), .B(OR4_289_Y), .C(OR4_169_Y), .D(
        OR4_220_Y), .Y(OR4_662_Y));
    OR4 OR4_439 (.A(OR4_15_Y), .B(OR4_267_Y), .C(OR4_566_Y), .D(
        OR4_134_Y), .Y(OR4_439_Y));
    OR4 OR4_346 (.A(\Z\R_DATA_TEMPR8[54] ), .B(\Z\R_DATA_TEMPR9[54] ), 
        .C(\Z\R_DATA_TEMPR10[54] ), .D(\Z\R_DATA_TEMPR11[54] ), .Y(
        OR4_346_Y));
    OR4 OR4_136 (.A(OR4_56_Y), .B(OR2_62_Y), .C(\Z\R_DATA_TEMPR22[4] ), 
        .D(\Z\R_DATA_TEMPR23[4] ), .Y(OR4_136_Y));
    OR2 OR2_20 (.A(\Z\R_DATA_TEMPR20[66] ), .B(\Z\R_DATA_TEMPR21[66] ), 
        .Y(OR2_20_Y));
    INV \INVBLKX1[0]  (.A(W_ADDR_c[10]), .Y(\Z\BLKX1[0] ));
    OR2 OR2_16 (.A(\Z\R_DATA_TEMPR20[48] ), .B(\Z\R_DATA_TEMPR21[48] ), 
        .Y(OR2_16_Y));
    CFG2 #( .INIT(4'h4) )  CFG2_6 (.A(R_ADDR_c[12]), .B(R_ADDR_c[11]), 
        .Y(CFG2_6_Y));
    OR2 OR2_27 (.A(\Z\R_DATA_TEMPR20[58] ), .B(\Z\R_DATA_TEMPR21[58] ), 
        .Y(OR2_27_Y));
    OR4 OR4_426 (.A(\Z\R_DATA_TEMPR0[67] ), .B(\Z\R_DATA_TEMPR1[67] ), 
        .C(\Z\R_DATA_TEMPR2[67] ), .D(\Z\R_DATA_TEMPR3[67] ), .Y(
        OR4_426_Y));
    CFG3 #( .INIT(8'h20) )  \CFG3_BLKY2[0]  (.A(CFG2_3_Y), .B(
        R_ADDR_c[13]), .C(R_EN_c), .Y(\Z\BLKY2[0] ));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%9%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0 (
        .A_DOUT({\Z\R_DATA_TEMPR9[39] , \Z\R_DATA_TEMPR9[38] , 
        \Z\R_DATA_TEMPR9[37] , \Z\R_DATA_TEMPR9[36] , 
        \Z\R_DATA_TEMPR9[35] , \Z\R_DATA_TEMPR9[34] , 
        \Z\R_DATA_TEMPR9[33] , \Z\R_DATA_TEMPR9[32] , 
        \Z\R_DATA_TEMPR9[31] , \Z\R_DATA_TEMPR9[30] , 
        \Z\R_DATA_TEMPR9[29] , \Z\R_DATA_TEMPR9[28] , 
        \Z\R_DATA_TEMPR9[27] , \Z\R_DATA_TEMPR9[26] , 
        \Z\R_DATA_TEMPR9[25] , \Z\R_DATA_TEMPR9[24] , 
        \Z\R_DATA_TEMPR9[23] , \Z\R_DATA_TEMPR9[22] , 
        \Z\R_DATA_TEMPR9[21] , \Z\R_DATA_TEMPR9[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR9[19] , \Z\R_DATA_TEMPR9[18] , 
        \Z\R_DATA_TEMPR9[17] , \Z\R_DATA_TEMPR9[16] , 
        \Z\R_DATA_TEMPR9[15] , \Z\R_DATA_TEMPR9[14] , 
        \Z\R_DATA_TEMPR9[13] , \Z\R_DATA_TEMPR9[12] , 
        \Z\R_DATA_TEMPR9[11] , \Z\R_DATA_TEMPR9[10] , 
        \Z\R_DATA_TEMPR9[9] , \Z\R_DATA_TEMPR9[8] , 
        \Z\R_DATA_TEMPR9[7] , \Z\R_DATA_TEMPR9[6] , 
        \Z\R_DATA_TEMPR9[5] , \Z\R_DATA_TEMPR9[4] , 
        \Z\R_DATA_TEMPR9[3] , \Z\R_DATA_TEMPR9[2] , 
        \Z\R_DATA_TEMPR9[1] , \Z\R_DATA_TEMPR9[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[9][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[2] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[2] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_203 (.A(\Z\R_DATA_TEMPR12[59] ), .B(\Z\R_DATA_TEMPR13[59] )
        , .C(\Z\R_DATA_TEMPR14[59] ), .D(\Z\R_DATA_TEMPR15[59] ), .Y(
        OR4_203_Y));
    OR4 OR4_290 (.A(\Z\R_DATA_TEMPR24[59] ), .B(\Z\R_DATA_TEMPR25[59] )
        , .C(\Z\R_DATA_TEMPR26[59] ), .D(\Z\R_DATA_TEMPR27[59] ), .Y(
        OR4_290_Y));
    OR4 OR4_597 (.A(\Z\R_DATA_TEMPR28[55] ), .B(\Z\R_DATA_TEMPR29[55] )
        , .C(\Z\R_DATA_TEMPR30[55] ), .D(\Z\R_DATA_TEMPR31[55] ), .Y(
        OR4_597_Y));
    OR4 OR4_338 (.A(OR4_111_Y), .B(OR4_694_Y), .C(OR4_574_Y), .D(
        OR4_609_Y), .Y(OR4_338_Y));
    OR4 OR4_273 (.A(\Z\R_DATA_TEMPR4[47] ), .B(\Z\R_DATA_TEMPR5[47] ), 
        .C(\Z\R_DATA_TEMPR6[47] ), .D(\Z\R_DATA_TEMPR7[47] ), .Y(
        OR4_273_Y));
    OR4 \OR4_R_DATA[77]  (.A(OR4_117_Y), .B(OR4_473_Y), .C(OR4_657_Y), 
        .D(OR4_717_Y), .Y(R_DATA_c[77]));
    OR4 OR4_322 (.A(\Z\R_DATA_TEMPR4[72] ), .B(\Z\R_DATA_TEMPR5[72] ), 
        .C(\Z\R_DATA_TEMPR6[72] ), .D(\Z\R_DATA_TEMPR7[72] ), .Y(
        OR4_322_Y));
    OR4 OR4_313 (.A(\Z\R_DATA_TEMPR4[18] ), .B(\Z\R_DATA_TEMPR5[18] ), 
        .C(\Z\R_DATA_TEMPR6[18] ), .D(\Z\R_DATA_TEMPR7[18] ), .Y(
        OR4_313_Y));
    OR4 OR4_710 (.A(\Z\R_DATA_TEMPR12[61] ), .B(\Z\R_DATA_TEMPR13[61] )
        , .C(\Z\R_DATA_TEMPR14[61] ), .D(\Z\R_DATA_TEMPR15[61] ), .Y(
        OR4_710_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%19%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0 (
        .A_DOUT({\Z\R_DATA_TEMPR19[39] , \Z\R_DATA_TEMPR19[38] , 
        \Z\R_DATA_TEMPR19[37] , \Z\R_DATA_TEMPR19[36] , 
        \Z\R_DATA_TEMPR19[35] , \Z\R_DATA_TEMPR19[34] , 
        \Z\R_DATA_TEMPR19[33] , \Z\R_DATA_TEMPR19[32] , 
        \Z\R_DATA_TEMPR19[31] , \Z\R_DATA_TEMPR19[30] , 
        \Z\R_DATA_TEMPR19[29] , \Z\R_DATA_TEMPR19[28] , 
        \Z\R_DATA_TEMPR19[27] , \Z\R_DATA_TEMPR19[26] , 
        \Z\R_DATA_TEMPR19[25] , \Z\R_DATA_TEMPR19[24] , 
        \Z\R_DATA_TEMPR19[23] , \Z\R_DATA_TEMPR19[22] , 
        \Z\R_DATA_TEMPR19[21] , \Z\R_DATA_TEMPR19[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR19[19] , \Z\R_DATA_TEMPR19[18] , 
        \Z\R_DATA_TEMPR19[17] , \Z\R_DATA_TEMPR19[16] , 
        \Z\R_DATA_TEMPR19[15] , \Z\R_DATA_TEMPR19[14] , 
        \Z\R_DATA_TEMPR19[13] , \Z\R_DATA_TEMPR19[12] , 
        \Z\R_DATA_TEMPR19[11] , \Z\R_DATA_TEMPR19[10] , 
        \Z\R_DATA_TEMPR19[9] , \Z\R_DATA_TEMPR19[8] , 
        \Z\R_DATA_TEMPR19[7] , \Z\R_DATA_TEMPR19[6] , 
        \Z\R_DATA_TEMPR19[5] , \Z\R_DATA_TEMPR19[4] , 
        \Z\R_DATA_TEMPR19[3] , \Z\R_DATA_TEMPR19[2] , 
        \Z\R_DATA_TEMPR19[1] , \Z\R_DATA_TEMPR19[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[19][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[4] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[4] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_699 (.A(\Z\R_DATA_TEMPR4[74] ), .B(\Z\R_DATA_TEMPR5[74] ), 
        .C(\Z\R_DATA_TEMPR6[74] ), .D(\Z\R_DATA_TEMPR7[74] ), .Y(
        OR4_699_Y));
    OR4 OR4_12 (.A(\Z\R_DATA_TEMPR0[58] ), .B(\Z\R_DATA_TEMPR1[58] ), 
        .C(\Z\R_DATA_TEMPR2[58] ), .D(\Z\R_DATA_TEMPR3[58] ), .Y(
        OR4_12_Y));
    OR4 OR4_583 (.A(\Z\R_DATA_TEMPR4[75] ), .B(\Z\R_DATA_TEMPR5[75] ), 
        .C(\Z\R_DATA_TEMPR6[75] ), .D(\Z\R_DATA_TEMPR7[75] ), .Y(
        OR4_583_Y));
    OR4 OR4_412 (.A(OR4_654_Y), .B(OR4_507_Y), .C(OR4_498_Y), .D(
        OR4_227_Y), .Y(OR4_412_Y));
    OR4 OR4_296 (.A(\Z\R_DATA_TEMPR12[49] ), .B(\Z\R_DATA_TEMPR13[49] )
        , .C(\Z\R_DATA_TEMPR14[49] ), .D(\Z\R_DATA_TEMPR15[49] ), .Y(
        OR4_296_Y));
    OR4 OR4_419 (.A(OR4_285_Y), .B(OR2_6_Y), .C(\Z\R_DATA_TEMPR22[33] )
        , .D(\Z\R_DATA_TEMPR23[33] ), .Y(OR4_419_Y));
    OR4 OR4_251 (.A(\Z\R_DATA_TEMPR16[55] ), .B(\Z\R_DATA_TEMPR17[55] )
        , .C(\Z\R_DATA_TEMPR18[55] ), .D(\Z\R_DATA_TEMPR19[55] ), .Y(
        OR4_251_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%11%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0 (
        .A_DOUT({\Z\R_DATA_TEMPR11[39] , \Z\R_DATA_TEMPR11[38] , 
        \Z\R_DATA_TEMPR11[37] , \Z\R_DATA_TEMPR11[36] , 
        \Z\R_DATA_TEMPR11[35] , \Z\R_DATA_TEMPR11[34] , 
        \Z\R_DATA_TEMPR11[33] , \Z\R_DATA_TEMPR11[32] , 
        \Z\R_DATA_TEMPR11[31] , \Z\R_DATA_TEMPR11[30] , 
        \Z\R_DATA_TEMPR11[29] , \Z\R_DATA_TEMPR11[28] , 
        \Z\R_DATA_TEMPR11[27] , \Z\R_DATA_TEMPR11[26] , 
        \Z\R_DATA_TEMPR11[25] , \Z\R_DATA_TEMPR11[24] , 
        \Z\R_DATA_TEMPR11[23] , \Z\R_DATA_TEMPR11[22] , 
        \Z\R_DATA_TEMPR11[21] , \Z\R_DATA_TEMPR11[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR11[19] , \Z\R_DATA_TEMPR11[18] , 
        \Z\R_DATA_TEMPR11[17] , \Z\R_DATA_TEMPR11[16] , 
        \Z\R_DATA_TEMPR11[15] , \Z\R_DATA_TEMPR11[14] , 
        \Z\R_DATA_TEMPR11[13] , \Z\R_DATA_TEMPR11[12] , 
        \Z\R_DATA_TEMPR11[11] , \Z\R_DATA_TEMPR11[10] , 
        \Z\R_DATA_TEMPR11[9] , \Z\R_DATA_TEMPR11[8] , 
        \Z\R_DATA_TEMPR11[7] , \Z\R_DATA_TEMPR11[6] , 
        \Z\R_DATA_TEMPR11[5] , \Z\R_DATA_TEMPR11[4] , 
        \Z\R_DATA_TEMPR11[3] , \Z\R_DATA_TEMPR11[2] , 
        \Z\R_DATA_TEMPR11[1] , \Z\R_DATA_TEMPR11[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[11][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[2] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[2] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_79 (.A(\Z\R_DATA_TEMPR8[50] ), .B(\Z\R_DATA_TEMPR9[50] ), 
        .C(\Z\R_DATA_TEMPR10[50] ), .D(\Z\R_DATA_TEMPR11[50] ), .Y(
        OR4_79_Y));
    OR4 OR4_139 (.A(\Z\R_DATA_TEMPR28[23] ), .B(\Z\R_DATA_TEMPR29[23] )
        , .C(\Z\R_DATA_TEMPR30[23] ), .D(\Z\R_DATA_TEMPR31[23] ), .Y(
        OR4_139_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%14%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C1 (
        .A_DOUT({\Z\R_DATA_TEMPR14[79] , \Z\R_DATA_TEMPR14[78] , 
        \Z\R_DATA_TEMPR14[77] , \Z\R_DATA_TEMPR14[76] , 
        \Z\R_DATA_TEMPR14[75] , \Z\R_DATA_TEMPR14[74] , 
        \Z\R_DATA_TEMPR14[73] , \Z\R_DATA_TEMPR14[72] , 
        \Z\R_DATA_TEMPR14[71] , \Z\R_DATA_TEMPR14[70] , 
        \Z\R_DATA_TEMPR14[69] , \Z\R_DATA_TEMPR14[68] , 
        \Z\R_DATA_TEMPR14[67] , \Z\R_DATA_TEMPR14[66] , 
        \Z\R_DATA_TEMPR14[65] , \Z\R_DATA_TEMPR14[64] , 
        \Z\R_DATA_TEMPR14[63] , \Z\R_DATA_TEMPR14[62] , 
        \Z\R_DATA_TEMPR14[61] , \Z\R_DATA_TEMPR14[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR14[59] , \Z\R_DATA_TEMPR14[58] , 
        \Z\R_DATA_TEMPR14[57] , \Z\R_DATA_TEMPR14[56] , 
        \Z\R_DATA_TEMPR14[55] , \Z\R_DATA_TEMPR14[54] , 
        \Z\R_DATA_TEMPR14[53] , \Z\R_DATA_TEMPR14[52] , 
        \Z\R_DATA_TEMPR14[51] , \Z\R_DATA_TEMPR14[50] , 
        \Z\R_DATA_TEMPR14[49] , \Z\R_DATA_TEMPR14[48] , 
        \Z\R_DATA_TEMPR14[47] , \Z\R_DATA_TEMPR14[46] , 
        \Z\R_DATA_TEMPR14[45] , \Z\R_DATA_TEMPR14[44] , 
        \Z\R_DATA_TEMPR14[43] , \Z\R_DATA_TEMPR14[42] , 
        \Z\R_DATA_TEMPR14[41] , \Z\R_DATA_TEMPR14[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[14][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[3] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[3] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_116 (.A(\Z\R_DATA_TEMPR0[33] ), .B(\Z\R_DATA_TEMPR1[33] ), 
        .C(\Z\R_DATA_TEMPR2[33] ), .D(\Z\R_DATA_TEMPR3[33] ), .Y(
        OR4_116_Y));
    OR4 OR4_608 (.A(OR4_245_Y), .B(OR4_17_Y), .C(OR4_52_Y), .D(
        OR4_192_Y), .Y(OR4_608_Y));
    OR4 OR4_144 (.A(\Z\R_DATA_TEMPR12[12] ), .B(\Z\R_DATA_TEMPR13[12] )
        , .C(\Z\R_DATA_TEMPR14[12] ), .D(\Z\R_DATA_TEMPR15[12] ), .Y(
        OR4_144_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%18%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0 (
        .A_DOUT({\Z\R_DATA_TEMPR18[39] , \Z\R_DATA_TEMPR18[38] , 
        \Z\R_DATA_TEMPR18[37] , \Z\R_DATA_TEMPR18[36] , 
        \Z\R_DATA_TEMPR18[35] , \Z\R_DATA_TEMPR18[34] , 
        \Z\R_DATA_TEMPR18[33] , \Z\R_DATA_TEMPR18[32] , 
        \Z\R_DATA_TEMPR18[31] , \Z\R_DATA_TEMPR18[30] , 
        \Z\R_DATA_TEMPR18[29] , \Z\R_DATA_TEMPR18[28] , 
        \Z\R_DATA_TEMPR18[27] , \Z\R_DATA_TEMPR18[26] , 
        \Z\R_DATA_TEMPR18[25] , \Z\R_DATA_TEMPR18[24] , 
        \Z\R_DATA_TEMPR18[23] , \Z\R_DATA_TEMPR18[22] , 
        \Z\R_DATA_TEMPR18[21] , \Z\R_DATA_TEMPR18[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR18[19] , \Z\R_DATA_TEMPR18[18] , 
        \Z\R_DATA_TEMPR18[17] , \Z\R_DATA_TEMPR18[16] , 
        \Z\R_DATA_TEMPR18[15] , \Z\R_DATA_TEMPR18[14] , 
        \Z\R_DATA_TEMPR18[13] , \Z\R_DATA_TEMPR18[12] , 
        \Z\R_DATA_TEMPR18[11] , \Z\R_DATA_TEMPR18[10] , 
        \Z\R_DATA_TEMPR18[9] , \Z\R_DATA_TEMPR18[8] , 
        \Z\R_DATA_TEMPR18[7] , \Z\R_DATA_TEMPR18[6] , 
        \Z\R_DATA_TEMPR18[5] , \Z\R_DATA_TEMPR18[4] , 
        \Z\R_DATA_TEMPR18[3] , \Z\R_DATA_TEMPR18[2] , 
        \Z\R_DATA_TEMPR18[1] , \Z\R_DATA_TEMPR18[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[18][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[4] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[4] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_694 (.A(\Z\R_DATA_TEMPR4[48] ), .B(\Z\R_DATA_TEMPR5[48] ), 
        .C(\Z\R_DATA_TEMPR6[48] ), .D(\Z\R_DATA_TEMPR7[48] ), .Y(
        OR4_694_Y));
    OR2 OR2_70 (.A(\Z\R_DATA_TEMPR20[43] ), .B(\Z\R_DATA_TEMPR21[43] ), 
        .Y(OR2_70_Y));
    OR4 OR4_678 (.A(\Z\R_DATA_TEMPR12[37] ), .B(\Z\R_DATA_TEMPR13[37] )
        , .C(\Z\R_DATA_TEMPR14[37] ), .D(\Z\R_DATA_TEMPR15[37] ), .Y(
        OR4_678_Y));
    OR4 OR4_602 (.A(\Z\R_DATA_TEMPR16[74] ), .B(\Z\R_DATA_TEMPR17[74] )
        , .C(\Z\R_DATA_TEMPR18[74] ), .D(\Z\R_DATA_TEMPR19[74] ), .Y(
        OR4_602_Y));
    OR4 \OR4_R_DATA[32]  (.A(OR4_690_Y), .B(OR4_672_Y), .C(OR4_567_Y), 
        .D(OR4_255_Y), .Y(R_DATA_c[32]));
    OR4 OR4_552 (.A(\Z\R_DATA_TEMPR4[25] ), .B(\Z\R_DATA_TEMPR5[25] ), 
        .C(\Z\R_DATA_TEMPR6[25] ), .D(\Z\R_DATA_TEMPR7[25] ), .Y(
        OR4_552_Y));
    OR2 OR2_77 (.A(\Z\R_DATA_TEMPR20[42] ), .B(\Z\R_DATA_TEMPR21[42] ), 
        .Y(OR2_77_Y));
    OR4 OR4_220 (.A(\Z\R_DATA_TEMPR12[78] ), .B(\Z\R_DATA_TEMPR13[78] )
        , .C(\Z\R_DATA_TEMPR14[78] ), .D(\Z\R_DATA_TEMPR15[78] ), .Y(
        OR4_220_Y));
    OR4 OR4_672 (.A(OR4_360_Y), .B(OR2_14_Y), .C(
        \Z\R_DATA_TEMPR22[32] ), .D(\Z\R_DATA_TEMPR23[32] ), .Y(
        OR4_672_Y));
    OR4 OR4_527 (.A(\Z\R_DATA_TEMPR4[32] ), .B(\Z\R_DATA_TEMPR5[32] ), 
        .C(\Z\R_DATA_TEMPR6[32] ), .D(\Z\R_DATA_TEMPR7[32] ), .Y(
        OR4_527_Y));
    OR4 OR4_318 (.A(\Z\R_DATA_TEMPR8[79] ), .B(\Z\R_DATA_TEMPR9[79] ), 
        .C(\Z\R_DATA_TEMPR10[79] ), .D(\Z\R_DATA_TEMPR11[79] ), .Y(
        OR4_318_Y));
    OR2 OR2_10 (.A(\Z\R_DATA_TEMPR20[9] ), .B(\Z\R_DATA_TEMPR21[9] ), 
        .Y(OR2_10_Y));
    OR4 \OR4_R_DATA[55]  (.A(OR4_181_Y), .B(OR4_520_Y), .C(OR4_70_Y), 
        .D(OR4_597_Y), .Y(R_DATA_c[55]));
    OR4 \OR4_R_DATA[3]  (.A(OR4_178_Y), .B(OR4_373_Y), .C(OR4_314_Y), 
        .D(OR4_371_Y), .Y(R_DATA_c[3]));
    OR2 OR2_17 (.A(\Z\R_DATA_TEMPR20[55] ), .B(\Z\R_DATA_TEMPR21[55] ), 
        .Y(OR2_17_Y));
    OR4 OR4_666 (.A(\Z\R_DATA_TEMPR4[24] ), .B(\Z\R_DATA_TEMPR5[24] ), 
        .C(\Z\R_DATA_TEMPR6[24] ), .D(\Z\R_DATA_TEMPR7[24] ), .Y(
        OR4_666_Y));
    OR4 OR4_629 (.A(\Z\R_DATA_TEMPR0[26] ), .B(\Z\R_DATA_TEMPR1[26] ), 
        .C(\Z\R_DATA_TEMPR2[26] ), .D(\Z\R_DATA_TEMPR3[26] ), .Y(
        OR4_629_Y));
    OR4 OR4_554 (.A(\Z\R_DATA_TEMPR4[27] ), .B(\Z\R_DATA_TEMPR5[27] ), 
        .C(\Z\R_DATA_TEMPR6[27] ), .D(\Z\R_DATA_TEMPR7[27] ), .Y(
        OR4_554_Y));
    OR4 OR4_546 (.A(\Z\R_DATA_TEMPR28[65] ), .B(\Z\R_DATA_TEMPR29[65] )
        , .C(\Z\R_DATA_TEMPR30[65] ), .D(\Z\R_DATA_TEMPR31[65] ), .Y(
        OR4_546_Y));
    OR4 OR4_226 (.A(\Z\R_DATA_TEMPR4[64] ), .B(\Z\R_DATA_TEMPR5[64] ), 
        .C(\Z\R_DATA_TEMPR6[64] ), .D(\Z\R_DATA_TEMPR7[64] ), .Y(
        OR4_226_Y));
    OR4 OR4_119 (.A(\Z\R_DATA_TEMPR24[37] ), .B(\Z\R_DATA_TEMPR25[37] )
        , .C(\Z\R_DATA_TEMPR26[37] ), .D(\Z\R_DATA_TEMPR27[37] ), .Y(
        OR4_119_Y));
    OR4 OR4_72 (.A(\Z\R_DATA_TEMPR0[50] ), .B(\Z\R_DATA_TEMPR1[50] ), 
        .C(\Z\R_DATA_TEMPR2[50] ), .D(\Z\R_DATA_TEMPR3[50] ), .Y(
        OR4_72_Y));
    OR4 OR4_637 (.A(\Z\R_DATA_TEMPR16[25] ), .B(\Z\R_DATA_TEMPR17[25] )
        , .C(\Z\R_DATA_TEMPR18[25] ), .D(\Z\R_DATA_TEMPR19[25] ), .Y(
        OR4_637_Y));
    OR4 OR4_624 (.A(\Z\R_DATA_TEMPR24[27] ), .B(\Z\R_DATA_TEMPR25[27] )
        , .C(\Z\R_DATA_TEMPR26[27] ), .D(\Z\R_DATA_TEMPR27[27] ), .Y(
        OR4_624_Y));
    OR4 OR4_351 (.A(\Z\R_DATA_TEMPR4[70] ), .B(\Z\R_DATA_TEMPR5[70] ), 
        .C(\Z\R_DATA_TEMPR6[70] ), .D(\Z\R_DATA_TEMPR7[70] ), .Y(
        OR4_351_Y));
    OR4 \OR4_R_DATA[33]  (.A(OR4_611_Y), .B(OR4_419_Y), .C(OR4_391_Y), 
        .D(OR4_366_Y), .Y(R_DATA_c[33]));
    OR2 OR2_28 (.A(\Z\R_DATA_TEMPR20[14] ), .B(\Z\R_DATA_TEMPR21[14] ), 
        .Y(OR2_28_Y));
    OR4 \OR4_R_DATA[25]  (.A(OR4_571_Y), .B(OR4_205_Y), .C(OR4_472_Y), 
        .D(OR4_274_Y), .Y(R_DATA_c[25]));
    OR4 OR4_450 (.A(\Z\R_DATA_TEMPR12[27] ), .B(\Z\R_DATA_TEMPR13[27] )
        , .C(\Z\R_DATA_TEMPR14[27] ), .D(\Z\R_DATA_TEMPR15[27] ), .Y(
        OR4_450_Y));
    OR4 OR4_283 (.A(\Z\R_DATA_TEMPR24[64] ), .B(\Z\R_DATA_TEMPR25[64] )
        , .C(\Z\R_DATA_TEMPR26[64] ), .D(\Z\R_DATA_TEMPR27[64] ), .Y(
        OR4_283_Y));
    OR4 OR4_96 (.A(\Z\R_DATA_TEMPR4[7] ), .B(\Z\R_DATA_TEMPR5[7] ), .C(
        \Z\R_DATA_TEMPR6[7] ), .D(\Z\R_DATA_TEMPR7[7] ), .Y(OR4_96_Y));
    OR4 OR4_548 (.A(\Z\R_DATA_TEMPR28[46] ), .B(\Z\R_DATA_TEMPR29[46] )
        , .C(\Z\R_DATA_TEMPR30[46] ), .D(\Z\R_DATA_TEMPR31[46] ), .Y(
        OR4_548_Y));
    OR4 OR4_54 (.A(\Z\R_DATA_TEMPR28[70] ), .B(\Z\R_DATA_TEMPR29[70] ), 
        .C(\Z\R_DATA_TEMPR30[70] ), .D(\Z\R_DATA_TEMPR31[70] ), .Y(
        OR4_54_Y));
    OR4 OR4_3 (.A(OR4_102_Y), .B(OR2_72_Y), .C(\Z\R_DATA_TEMPR22[70] ), 
        .D(\Z\R_DATA_TEMPR23[70] ), .Y(OR4_3_Y));
    OR4 OR4_364 (.A(\Z\R_DATA_TEMPR12[60] ), .B(\Z\R_DATA_TEMPR13[60] )
        , .C(\Z\R_DATA_TEMPR14[60] ), .D(\Z\R_DATA_TEMPR15[60] ), .Y(
        OR4_364_Y));
    OR4 OR4_606 (.A(\Z\R_DATA_TEMPR16[69] ), .B(\Z\R_DATA_TEMPR17[69] )
        , .C(\Z\R_DATA_TEMPR18[69] ), .D(\Z\R_DATA_TEMPR19[69] ), .Y(
        OR4_606_Y));
    OR4 OR4_715 (.A(OR4_616_Y), .B(OR2_78_Y), .C(
        \Z\R_DATA_TEMPR22[67] ), .D(\Z\R_DATA_TEMPR23[67] ), .Y(
        OR4_715_Y));
    OR4 OR4_617 (.A(\Z\R_DATA_TEMPR12[79] ), .B(\Z\R_DATA_TEMPR13[79] )
        , .C(\Z\R_DATA_TEMPR14[79] ), .D(\Z\R_DATA_TEMPR15[79] ), .Y(
        OR4_617_Y));
    OR4 OR4_446 (.A(\Z\R_DATA_TEMPR8[26] ), .B(\Z\R_DATA_TEMPR9[26] ), 
        .C(\Z\R_DATA_TEMPR10[26] ), .D(\Z\R_DATA_TEMPR11[26] ), .Y(
        OR4_446_Y));
    OR4 OR4_161 (.A(\Z\R_DATA_TEMPR0[75] ), .B(\Z\R_DATA_TEMPR1[75] ), 
        .C(\Z\R_DATA_TEMPR2[75] ), .D(\Z\R_DATA_TEMPR3[75] ), .Y(
        OR4_161_Y));
    OR4 OR4_716 (.A(OR4_408_Y), .B(OR2_41_Y), .C(
        \Z\R_DATA_TEMPR22[62] ), .D(\Z\R_DATA_TEMPR23[62] ), .Y(
        OR4_716_Y));
    OR4 OR4_676 (.A(\Z\R_DATA_TEMPR8[36] ), .B(\Z\R_DATA_TEMPR9[36] ), 
        .C(\Z\R_DATA_TEMPR10[36] ), .D(\Z\R_DATA_TEMPR11[36] ), .Y(
        OR4_676_Y));
    OR4 OR4_237 (.A(\Z\R_DATA_TEMPR12[25] ), .B(\Z\R_DATA_TEMPR13[25] )
        , .C(\Z\R_DATA_TEMPR14[25] ), .D(\Z\R_DATA_TEMPR15[25] ), .Y(
        OR4_237_Y));
    OR4 OR4_688 (.A(OR4_105_Y), .B(OR2_13_Y), .C(\Z\R_DATA_TEMPR22[5] )
        , .D(\Z\R_DATA_TEMPR23[5] ), .Y(OR4_688_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%23%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0 (
        .A_DOUT({\Z\R_DATA_TEMPR23[39] , \Z\R_DATA_TEMPR23[38] , 
        \Z\R_DATA_TEMPR23[37] , \Z\R_DATA_TEMPR23[36] , 
        \Z\R_DATA_TEMPR23[35] , \Z\R_DATA_TEMPR23[34] , 
        \Z\R_DATA_TEMPR23[33] , \Z\R_DATA_TEMPR23[32] , 
        \Z\R_DATA_TEMPR23[31] , \Z\R_DATA_TEMPR23[30] , 
        \Z\R_DATA_TEMPR23[29] , \Z\R_DATA_TEMPR23[28] , 
        \Z\R_DATA_TEMPR23[27] , \Z\R_DATA_TEMPR23[26] , 
        \Z\R_DATA_TEMPR23[25] , \Z\R_DATA_TEMPR23[24] , 
        \Z\R_DATA_TEMPR23[23] , \Z\R_DATA_TEMPR23[22] , 
        \Z\R_DATA_TEMPR23[21] , \Z\R_DATA_TEMPR23[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR23[19] , \Z\R_DATA_TEMPR23[18] , 
        \Z\R_DATA_TEMPR23[17] , \Z\R_DATA_TEMPR23[16] , 
        \Z\R_DATA_TEMPR23[15] , \Z\R_DATA_TEMPR23[14] , 
        \Z\R_DATA_TEMPR23[13] , \Z\R_DATA_TEMPR23[12] , 
        \Z\R_DATA_TEMPR23[11] , \Z\R_DATA_TEMPR23[10] , 
        \Z\R_DATA_TEMPR23[9] , \Z\R_DATA_TEMPR23[8] , 
        \Z\R_DATA_TEMPR23[7] , \Z\R_DATA_TEMPR23[6] , 
        \Z\R_DATA_TEMPR23[5] , \Z\R_DATA_TEMPR23[4] , 
        \Z\R_DATA_TEMPR23[3] , \Z\R_DATA_TEMPR23[2] , 
        \Z\R_DATA_TEMPR23[1] , \Z\R_DATA_TEMPR23[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[23][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[5] , R_ADDR_c[10], 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[5] , W_ADDR_c[10], 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_137 (.A(\Z\R_DATA_TEMPR8[77] ), .B(\Z\R_DATA_TEMPR9[77] ), 
        .C(\Z\R_DATA_TEMPR10[77] ), .D(\Z\R_DATA_TEMPR11[77] ), .Y(
        OR4_137_Y));
    OR2 OR2_78 (.A(\Z\R_DATA_TEMPR20[67] ), .B(\Z\R_DATA_TEMPR21[67] ), 
        .Y(OR2_78_Y));
    OR4 OR4_682 (.A(\Z\R_DATA_TEMPR24[17] ), .B(\Z\R_DATA_TEMPR25[17] )
        , .C(\Z\R_DATA_TEMPR26[17] ), .D(\Z\R_DATA_TEMPR27[17] ), .Y(
        OR4_682_Y));
    OR4 OR4_342 (.A(\Z\R_DATA_TEMPR4[71] ), .B(\Z\R_DATA_TEMPR5[71] ), 
        .C(\Z\R_DATA_TEMPR6[71] ), .D(\Z\R_DATA_TEMPR7[71] ), .Y(
        OR4_342_Y));
    OR4 OR4_461 (.A(\Z\R_DATA_TEMPR16[52] ), .B(\Z\R_DATA_TEMPR17[52] )
        , .C(\Z\R_DATA_TEMPR18[52] ), .D(\Z\R_DATA_TEMPR19[52] ), .Y(
        OR4_461_Y));
    OR4 OR4_359 (.A(\Z\R_DATA_TEMPR24[10] ), .B(\Z\R_DATA_TEMPR25[10] )
        , .C(\Z\R_DATA_TEMPR26[10] ), .D(\Z\R_DATA_TEMPR27[10] ), .Y(
        OR4_359_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%6%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C1 (
        .A_DOUT({\Z\R_DATA_TEMPR6[79] , \Z\R_DATA_TEMPR6[78] , 
        \Z\R_DATA_TEMPR6[77] , \Z\R_DATA_TEMPR6[76] , 
        \Z\R_DATA_TEMPR6[75] , \Z\R_DATA_TEMPR6[74] , 
        \Z\R_DATA_TEMPR6[73] , \Z\R_DATA_TEMPR6[72] , 
        \Z\R_DATA_TEMPR6[71] , \Z\R_DATA_TEMPR6[70] , 
        \Z\R_DATA_TEMPR6[69] , \Z\R_DATA_TEMPR6[68] , 
        \Z\R_DATA_TEMPR6[67] , \Z\R_DATA_TEMPR6[66] , 
        \Z\R_DATA_TEMPR6[65] , \Z\R_DATA_TEMPR6[64] , 
        \Z\R_DATA_TEMPR6[63] , \Z\R_DATA_TEMPR6[62] , 
        \Z\R_DATA_TEMPR6[61] , \Z\R_DATA_TEMPR6[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR6[59] , \Z\R_DATA_TEMPR6[58] , 
        \Z\R_DATA_TEMPR6[57] , \Z\R_DATA_TEMPR6[56] , 
        \Z\R_DATA_TEMPR6[55] , \Z\R_DATA_TEMPR6[54] , 
        \Z\R_DATA_TEMPR6[53] , \Z\R_DATA_TEMPR6[52] , 
        \Z\R_DATA_TEMPR6[51] , \Z\R_DATA_TEMPR6[50] , 
        \Z\R_DATA_TEMPR6[49] , \Z\R_DATA_TEMPR6[48] , 
        \Z\R_DATA_TEMPR6[47] , \Z\R_DATA_TEMPR6[46] , 
        \Z\R_DATA_TEMPR6[45] , \Z\R_DATA_TEMPR6[44] , 
        \Z\R_DATA_TEMPR6[43] , \Z\R_DATA_TEMPR6[42] , 
        \Z\R_DATA_TEMPR6[41] , \Z\R_DATA_TEMPR6[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[6][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[1] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[1] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_14 (.A(\Z\R_DATA_TEMPR0[34] ), .B(\Z\R_DATA_TEMPR1[34] ), 
        .C(\Z\R_DATA_TEMPR2[34] ), .D(\Z\R_DATA_TEMPR3[34] ), .Y(
        OR4_14_Y));
    OR4 OR4_468 (.A(OR4_198_Y), .B(OR2_53_Y), .C(
        \Z\R_DATA_TEMPR22[65] ), .D(\Z\R_DATA_TEMPR23[65] ), .Y(
        OR4_468_Y));
    OR2 OR2_18 (.A(\Z\R_DATA_TEMPR20[15] ), .B(\Z\R_DATA_TEMPR21[15] ), 
        .Y(OR2_18_Y));
    OR4 OR4_291 (.A(\Z\R_DATA_TEMPR8[45] ), .B(\Z\R_DATA_TEMPR9[45] ), 
        .C(\Z\R_DATA_TEMPR10[45] ), .D(\Z\R_DATA_TEMPR11[45] ), .Y(
        OR4_291_Y));
    OR4 OR4_234 (.A(OR4_667_Y), .B(OR2_73_Y), .C(
        \Z\R_DATA_TEMPR22[75] ), .D(\Z\R_DATA_TEMPR23[75] ), .Y(
        OR4_234_Y));
    OR4 OR4_90 (.A(OR4_239_Y), .B(OR4_639_Y), .C(OR4_399_Y), .D(
        OR4_157_Y), .Y(OR4_90_Y));
    OR4 OR4_46 (.A(\Z\R_DATA_TEMPR16[47] ), .B(\Z\R_DATA_TEMPR17[47] ), 
        .C(\Z\R_DATA_TEMPR18[47] ), .D(\Z\R_DATA_TEMPR19[47] ), .Y(
        OR4_46_Y));
    OR4 OR4_97 (.A(\Z\R_DATA_TEMPR24[76] ), .B(\Z\R_DATA_TEMPR25[76] ), 
        .C(\Z\R_DATA_TEMPR26[76] ), .D(\Z\R_DATA_TEMPR27[76] ), .Y(
        OR4_97_Y));
    OR4 OR4_569 (.A(\Z\R_DATA_TEMPR16[24] ), .B(\Z\R_DATA_TEMPR17[24] )
        , .C(\Z\R_DATA_TEMPR18[24] ), .D(\Z\R_DATA_TEMPR19[24] ), .Y(
        OR4_569_Y));
    OR4 \OR4_R_DATA[6]  (.A(OR4_168_Y), .B(OR4_515_Y), .C(OR4_27_Y), 
        .D(OR4_118_Y), .Y(R_DATA_c[6]));
    OR4 OR4_63 (.A(\Z\R_DATA_TEMPR8[1] ), .B(\Z\R_DATA_TEMPR9[1] ), .C(
        \Z\R_DATA_TEMPR10[1] ), .D(\Z\R_DATA_TEMPR11[1] ), .Y(OR4_63_Y)
        );
    OR4 OR4_592 (.A(\Z\R_DATA_TEMPR28[0] ), .B(\Z\R_DATA_TEMPR29[0] ), 
        .C(\Z\R_DATA_TEMPR30[0] ), .D(\Z\R_DATA_TEMPR31[0] ), .Y(
        OR4_592_Y));
    OR4 OR4_560 (.A(\Z\R_DATA_TEMPR28[9] ), .B(\Z\R_DATA_TEMPR29[9] ), 
        .C(\Z\R_DATA_TEMPR30[9] ), .D(\Z\R_DATA_TEMPR31[9] ), .Y(
        OR4_560_Y));
    OR4 OR4_217 (.A(\Z\R_DATA_TEMPR24[28] ), .B(\Z\R_DATA_TEMPR25[28] )
        , .C(\Z\R_DATA_TEMPR26[28] ), .D(\Z\R_DATA_TEMPR27[28] ), .Y(
        OR4_217_Y));
    OR4 OR4_304 (.A(\Z\R_DATA_TEMPR4[59] ), .B(\Z\R_DATA_TEMPR5[59] ), 
        .C(\Z\R_DATA_TEMPR6[59] ), .D(\Z\R_DATA_TEMPR7[59] ), .Y(
        OR4_304_Y));
    OR4 OR4_240 (.A(OR4_524_Y), .B(OR4_40_Y), .C(OR4_347_Y), .D(
        OR4_649_Y), .Y(OR4_240_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%20%1%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C1 (
        .A_DOUT({\Z\R_DATA_TEMPR20[79] , \Z\R_DATA_TEMPR20[78] , 
        \Z\R_DATA_TEMPR20[77] , \Z\R_DATA_TEMPR20[76] , 
        \Z\R_DATA_TEMPR20[75] , \Z\R_DATA_TEMPR20[74] , 
        \Z\R_DATA_TEMPR20[73] , \Z\R_DATA_TEMPR20[72] , 
        \Z\R_DATA_TEMPR20[71] , \Z\R_DATA_TEMPR20[70] , 
        \Z\R_DATA_TEMPR20[69] , \Z\R_DATA_TEMPR20[68] , 
        \Z\R_DATA_TEMPR20[67] , \Z\R_DATA_TEMPR20[66] , 
        \Z\R_DATA_TEMPR20[65] , \Z\R_DATA_TEMPR20[64] , 
        \Z\R_DATA_TEMPR20[63] , \Z\R_DATA_TEMPR20[62] , 
        \Z\R_DATA_TEMPR20[61] , \Z\R_DATA_TEMPR20[60] }), .B_DOUT({
        \Z\R_DATA_TEMPR20[59] , \Z\R_DATA_TEMPR20[58] , 
        \Z\R_DATA_TEMPR20[57] , \Z\R_DATA_TEMPR20[56] , 
        \Z\R_DATA_TEMPR20[55] , \Z\R_DATA_TEMPR20[54] , 
        \Z\R_DATA_TEMPR20[53] , \Z\R_DATA_TEMPR20[52] , 
        \Z\R_DATA_TEMPR20[51] , \Z\R_DATA_TEMPR20[50] , 
        \Z\R_DATA_TEMPR20[49] , \Z\R_DATA_TEMPR20[48] , 
        \Z\R_DATA_TEMPR20[47] , \Z\R_DATA_TEMPR20[46] , 
        \Z\R_DATA_TEMPR20[45] , \Z\R_DATA_TEMPR20[44] , 
        \Z\R_DATA_TEMPR20[43] , \Z\R_DATA_TEMPR20[42] , 
        \Z\R_DATA_TEMPR20[41] , \Z\R_DATA_TEMPR20[40] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C1_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C1_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[20][1] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[5] , \Z\BLKY1[0] , 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[79], 
        W_DATA_c[78], W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], 
        W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], 
        W_DATA_c[70], W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[7], WBYTE_EN_c[6]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[5] , \Z\BLKX1[0] , 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[59], 
        W_DATA_c[58], W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], 
        W_DATA_c[54], W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], 
        W_DATA_c[50], W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], 
        W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], 
        W_DATA_c[42], W_DATA_c[41], W_DATA_c[40]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN_c[5], WBYTE_EN_c[4]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_117 (.A(OR4_195_Y), .B(OR4_584_Y), .C(OR4_137_Y), .D(
        OR4_489_Y), .Y(OR4_117_Y));
    OR4 OR4_547 (.A(\Z\R_DATA_TEMPR28[34] ), .B(\Z\R_DATA_TEMPR29[34] )
        , .C(\Z\R_DATA_TEMPR30[34] ), .D(\Z\R_DATA_TEMPR31[34] ), .Y(
        OR4_547_Y));
    OR4 OR4_335 (.A(OR4_232_Y), .B(OR4_376_Y), .C(OR4_451_Y), .D(
        OR4_270_Y), .Y(OR4_335_Y));
    OR4 \OR4_R_DATA[1]  (.A(OR4_589_Y), .B(OR4_677_Y), .C(OR4_480_Y), 
        .D(OR4_384_Y), .Y(R_DATA_c[1]));
    OR4 OR4_374 (.A(OR4_569_Y), .B(OR2_51_Y), .C(
        \Z\R_DATA_TEMPR22[24] ), .D(\Z\R_DATA_TEMPR23[24] ), .Y(
        OR4_374_Y));
    OR4 OR4_101 (.A(\Z\R_DATA_TEMPR28[26] ), .B(\Z\R_DATA_TEMPR29[26] )
        , .C(\Z\R_DATA_TEMPR30[26] ), .D(\Z\R_DATA_TEMPR31[26] ), .Y(
        OR4_101_Y));
    OR4 OR4_649 (.A(\Z\R_DATA_TEMPR12[19] ), .B(\Z\R_DATA_TEMPR13[19] )
        , .C(\Z\R_DATA_TEMPR14[19] ), .D(\Z\R_DATA_TEMPR15[19] ), .Y(
        OR4_649_Y));
    OR4 OR4_594 (.A(OR4_222_Y), .B(OR2_29_Y), .C(
        \Z\R_DATA_TEMPR22[18] ), .D(\Z\R_DATA_TEMPR23[18] ), .Y(
        OR4_594_Y));
    OR4 OR4_171 (.A(OR4_458_Y), .B(OR4_704_Y), .C(OR4_288_Y), .D(
        OR4_585_Y), .Y(OR4_171_Y));
    OR4 OR4_713 (.A(OR4_334_Y), .B(OR4_114_Y), .C(OR4_160_Y), .D(
        OR4_287_Y), .Y(OR4_713_Y));
    OR4 OR4_553 (.A(\Z\R_DATA_TEMPR16[46] ), .B(\Z\R_DATA_TEMPR17[46] )
        , .C(\Z\R_DATA_TEMPR18[46] ), .D(\Z\R_DATA_TEMPR19[46] ), .Y(
        OR4_553_Y));
    OR4 OR4_214 (.A(OR4_306_Y), .B(OR2_25_Y), .C(
        \Z\R_DATA_TEMPR22[30] ), .D(\Z\R_DATA_TEMPR23[30] ), .Y(
        OR4_214_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%10%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0 (
        .A_DOUT({\Z\R_DATA_TEMPR10[39] , \Z\R_DATA_TEMPR10[38] , 
        \Z\R_DATA_TEMPR10[37] , \Z\R_DATA_TEMPR10[36] , 
        \Z\R_DATA_TEMPR10[35] , \Z\R_DATA_TEMPR10[34] , 
        \Z\R_DATA_TEMPR10[33] , \Z\R_DATA_TEMPR10[32] , 
        \Z\R_DATA_TEMPR10[31] , \Z\R_DATA_TEMPR10[30] , 
        \Z\R_DATA_TEMPR10[29] , \Z\R_DATA_TEMPR10[28] , 
        \Z\R_DATA_TEMPR10[27] , \Z\R_DATA_TEMPR10[26] , 
        \Z\R_DATA_TEMPR10[25] , \Z\R_DATA_TEMPR10[24] , 
        \Z\R_DATA_TEMPR10[23] , \Z\R_DATA_TEMPR10[22] , 
        \Z\R_DATA_TEMPR10[21] , \Z\R_DATA_TEMPR10[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR10[19] , \Z\R_DATA_TEMPR10[18] , 
        \Z\R_DATA_TEMPR10[17] , \Z\R_DATA_TEMPR10[16] , 
        \Z\R_DATA_TEMPR10[15] , \Z\R_DATA_TEMPR10[14] , 
        \Z\R_DATA_TEMPR10[13] , \Z\R_DATA_TEMPR10[12] , 
        \Z\R_DATA_TEMPR10[11] , \Z\R_DATA_TEMPR10[10] , 
        \Z\R_DATA_TEMPR10[9] , \Z\R_DATA_TEMPR10[8] , 
        \Z\R_DATA_TEMPR10[7] , \Z\R_DATA_TEMPR10[6] , 
        \Z\R_DATA_TEMPR10[5] , \Z\R_DATA_TEMPR10[4] , 
        \Z\R_DATA_TEMPR10[3] , \Z\R_DATA_TEMPR10[2] , 
        \Z\R_DATA_TEMPR10[1] , \Z\R_DATA_TEMPR10[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[10][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[2] , R_ADDR_c[10], 
        \Z\BLKY0[0] }), .A_CLK(CLK), .A_DIN({W_DATA_c[39], 
        W_DATA_c[38], W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], 
        W_DATA_c[34], W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], 
        W_DATA_c[30], W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], 
        W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], 
        W_DATA_c[22], W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), 
        .A_WEN({WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[2] , W_ADDR_c[10], 
        \Z\BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA_c[19], 
        W_DATA_c[18], W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], 
        W_DATA_c[14], W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], 
        W_DATA_c[10], W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], 
        W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], 
        W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({
        WBYTE_EN_c[1], WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(GND), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(GND), .ECC_BYPASS(GND));
    OR4 OR4_246 (.A(\Z\R_DATA_TEMPR24[4] ), .B(\Z\R_DATA_TEMPR25[4] ), 
        .C(\Z\R_DATA_TEMPR26[4] ), .D(\Z\R_DATA_TEMPR27[4] ), .Y(
        OR4_246_Y));
    OR4 OR4_221 (.A(\Z\R_DATA_TEMPR4[39] ), .B(\Z\R_DATA_TEMPR5[39] ), 
        .C(\Z\R_DATA_TEMPR6[39] ), .D(\Z\R_DATA_TEMPR7[39] ), .Y(
        OR4_221_Y));
    OR4 OR4_401 (.A(\Z\R_DATA_TEMPR24[56] ), .B(\Z\R_DATA_TEMPR25[56] )
        , .C(\Z\R_DATA_TEMPR26[56] ), .D(\Z\R_DATA_TEMPR27[56] ), .Y(
        OR4_401_Y));
    OR4 \OR4_R_DATA[58]  (.A(OR4_249_Y), .B(OR4_133_Y), .C(OR4_532_Y), 
        .D(OR4_634_Y), .Y(R_DATA_c[58]));
    OR4 OR4_74 (.A(\Z\R_DATA_TEMPR16[20] ), .B(\Z\R_DATA_TEMPR17[20] ), 
        .C(\Z\R_DATA_TEMPR18[20] ), .D(\Z\R_DATA_TEMPR19[20] ), .Y(
        OR4_74_Y));
    OR4 OR4_408 (.A(\Z\R_DATA_TEMPR16[62] ), .B(\Z\R_DATA_TEMPR17[62] )
        , .C(\Z\R_DATA_TEMPR18[62] ), .D(\Z\R_DATA_TEMPR19[62] ), .Y(
        OR4_408_Y));
    CFG3 #( .INIT(8'h80) )  \CFG3_BLKX2[6]  (.A(CFG2_7_Y), .B(
        W_ADDR_c[13]), .C(W_EN_c), .Y(\Z\BLKX2[6] ));
    OR4 OR4_471 (.A(\Z\R_DATA_TEMPR4[16] ), .B(\Z\R_DATA_TEMPR5[16] ), 
        .C(\Z\R_DATA_TEMPR6[16] ), .D(\Z\R_DATA_TEMPR7[16] ), .Y(
        OR4_471_Y));
    OR4 OR4_363 (.A(\Z\R_DATA_TEMPR12[62] ), .B(\Z\R_DATA_TEMPR13[62] )
        , .C(\Z\R_DATA_TEMPR14[62] ), .D(\Z\R_DATA_TEMPR15[62] ), .Y(
        OR4_363_Y));
    OR4 OR4_478 (.A(\Z\R_DATA_TEMPR8[2] ), .B(\Z\R_DATA_TEMPR9[2] ), 
        .C(\Z\R_DATA_TEMPR10[2] ), .D(\Z\R_DATA_TEMPR11[2] ), .Y(
        OR4_478_Y));
    OR4 OR4_391 (.A(\Z\R_DATA_TEMPR24[33] ), .B(\Z\R_DATA_TEMPR25[33] )
        , .C(\Z\R_DATA_TEMPR26[33] ), .D(\Z\R_DATA_TEMPR27[33] ), .Y(
        OR4_391_Y));
    OR4 OR4_644 (.A(\Z\R_DATA_TEMPR4[36] ), .B(\Z\R_DATA_TEMPR5[36] ), 
        .C(\Z\R_DATA_TEMPR6[36] ), .D(\Z\R_DATA_TEMPR7[36] ), .Y(
        OR4_644_Y));
    OR4 OR4_61 (.A(\Z\R_DATA_TEMPR0[59] ), .B(\Z\R_DATA_TEMPR1[59] ), 
        .C(\Z\R_DATA_TEMPR2[59] ), .D(\Z\R_DATA_TEMPR3[59] ), .Y(
        OR4_61_Y));
    OR4 OR4_462 (.A(OR4_596_Y), .B(OR4_297_Y), .C(OR4_445_Y), .D(
        OR4_80_Y), .Y(OR4_462_Y));
    OR4 OR4_635 (.A(OR4_110_Y), .B(OR2_56_Y), .C(
        \Z\R_DATA_TEMPR22[21] ), .D(\Z\R_DATA_TEMPR23[21] ), .Y(
        OR4_635_Y));
    OR4 OR4_522 (.A(\Z\R_DATA_TEMPR12[42] ), .B(\Z\R_DATA_TEMPR13[42] )
        , .C(\Z\R_DATA_TEMPR14[42] ), .D(\Z\R_DATA_TEMPR15[42] ), .Y(
        OR4_522_Y));
    OR4 OR4_686 (.A(OR4_572_Y), .B(OR4_718_Y), .C(OR4_71_Y), .D(
        OR4_610_Y), .Y(OR4_686_Y));
    OR4 OR4_469 (.A(OR4_333_Y), .B(OR2_34_Y), .C(
        \Z\R_DATA_TEMPR22[63] ), .D(\Z\R_DATA_TEMPR23[63] ), .Y(
        OR4_469_Y));
    OR4 OR4_315 (.A(\Z\R_DATA_TEMPR28[24] ), .B(\Z\R_DATA_TEMPR29[24] )
        , .C(\Z\R_DATA_TEMPR30[24] ), .D(\Z\R_DATA_TEMPR31[24] ), .Y(
        OR4_315_Y));
    OR2 OR2_5 (.A(\Z\R_DATA_TEMPR20[40] ), .B(\Z\R_DATA_TEMPR21[40] ), 
        .Y(OR2_5_Y));
    OR4 OR4_490 (.A(\Z\R_DATA_TEMPR16[2] ), .B(\Z\R_DATA_TEMPR17[2] ), 
        .C(\Z\R_DATA_TEMPR18[2] ), .D(\Z\R_DATA_TEMPR19[2] ), .Y(
        OR4_490_Y));
    OR4 OR4_40 (.A(\Z\R_DATA_TEMPR4[19] ), .B(\Z\R_DATA_TEMPR5[19] ), 
        .C(\Z\R_DATA_TEMPR6[19] ), .D(\Z\R_DATA_TEMPR7[19] ), .Y(
        OR4_40_Y));
    RAM1K20 #( .MEMORYFILE(""), .RAMINDEX("PF_SRAM_AHBL_AXI_C1%16384-16384%80-80%POWER%5%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0 (
        .A_DOUT({\Z\R_DATA_TEMPR5[39] , \Z\R_DATA_TEMPR5[38] , 
        \Z\R_DATA_TEMPR5[37] , \Z\R_DATA_TEMPR5[36] , 
        \Z\R_DATA_TEMPR5[35] , \Z\R_DATA_TEMPR5[34] , 
        \Z\R_DATA_TEMPR5[33] , \Z\R_DATA_TEMPR5[32] , 
        \Z\R_DATA_TEMPR5[31] , \Z\R_DATA_TEMPR5[30] , 
        \Z\R_DATA_TEMPR5[29] , \Z\R_DATA_TEMPR5[28] , 
        \Z\R_DATA_TEMPR5[27] , \Z\R_DATA_TEMPR5[26] , 
        \Z\R_DATA_TEMPR5[25] , \Z\R_DATA_TEMPR5[24] , 
        \Z\R_DATA_TEMPR5[23] , \Z\R_DATA_TEMPR5[22] , 
        \Z\R_DATA_TEMPR5[21] , \Z\R_DATA_TEMPR5[20] }), .B_DOUT({
        \Z\R_DATA_TEMPR5[19] , \Z\R_DATA_TEMPR5[18] , 
        \Z\R_DATA_TEMPR5[17] , \Z\R_DATA_TEMPR5[16] , 
        \Z\R_DATA_TEMPR5[15] , \Z\R_DATA_TEMPR5[14] , 
        \Z\R_DATA_TEMPR5[13] , \Z\R_DATA_TEMPR5[12] , 
        \Z\R_DATA_TEMPR5[11] , \Z\R_DATA_TEMPR5[10] , 
        \Z\R_DATA_TEMPR5[9] , \Z\R_DATA_TEMPR5[8] , 
        \Z\R_DATA_TEMPR5[7] , \Z\R_DATA_TEMPR5[6] , 
        \Z\R_DATA_TEMPR5[5] , \Z\R_DATA_TEMPR5[4] , 
        \Z\R_DATA_TEMPR5[3] , \Z\R_DATA_TEMPR5[2] , 
        \Z\R_DATA_TEMPR5[1] , \Z\R_DATA_TEMPR5[0] }), .DB_DETECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0_DB_DETECT)
        , .SB_CORRECT(
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0_SB_CORRECT)
        , .ACCESS_BUSY(\Z\ACCESS_BUSY[5][0] ), .A_ADDR({R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .A_BLK_EN({\Z\BLKY2[1] , \Z\BLKY1[0] , 
        R_ADDR_c[9]}), .A_CLK(CLK), .A_DIN({W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20]}), .A_REN(VCC), .A_WEN({
        WBYTE_EN_c[3], WBYTE_EN_c[2]}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR_c[8], 
        W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], 
        W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0], GND, GND, 
        GND, GND, GND}), .B_BLK_EN({\Z\BLKX2[1] , \Z\BLKX1[0] , 
        W_ADDR_c[9]}), .B_CLK(CLK), .B_DIN({W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(GND), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(GND)
        , .ECC_BYPASS(GND));
    OR4 OR4_509 (.A(\Z\R_DATA_TEMPR8[16] ), .B(\Z\R_DATA_TEMPR9[16] ), 
        .C(\Z\R_DATA_TEMPR10[16] ), .D(\Z\R_DATA_TEMPR11[16] ), .Y(
        OR4_509_Y));
    OR4 OR4_166 (.A(\Z\R_DATA_TEMPR4[34] ), .B(\Z\R_DATA_TEMPR5[34] ), 
        .C(\Z\R_DATA_TEMPR6[34] ), .D(\Z\R_DATA_TEMPR7[34] ), .Y(
        OR4_166_Y));
    OR4 OR4_500 (.A(\Z\R_DATA_TEMPR12[58] ), .B(\Z\R_DATA_TEMPR13[58] )
        , .C(\Z\R_DATA_TEMPR14[58] ), .D(\Z\R_DATA_TEMPR15[58] ), .Y(
        OR4_500_Y));
    OR4 OR4_47 (.A(\Z\R_DATA_TEMPR12[34] ), .B(\Z\R_DATA_TEMPR13[34] ), 
        .C(\Z\R_DATA_TEMPR14[34] ), .D(\Z\R_DATA_TEMPR15[34] ), .Y(
        OR4_47_Y));
    OR4 OR4_579 (.A(\Z\R_DATA_TEMPR12[26] ), .B(\Z\R_DATA_TEMPR13[26] )
        , .C(\Z\R_DATA_TEMPR14[26] ), .D(\Z\R_DATA_TEMPR15[26] ), .Y(
        OR4_579_Y));
    OR4 OR4_570 (.A(\Z\R_DATA_TEMPR16[42] ), .B(\Z\R_DATA_TEMPR17[42] )
        , .C(\Z\R_DATA_TEMPR18[42] ), .D(\Z\R_DATA_TEMPR19[42] ), .Y(
        OR4_570_Y));
    OR4 OR4_524 (.A(\Z\R_DATA_TEMPR0[19] ), .B(\Z\R_DATA_TEMPR1[19] ), 
        .C(\Z\R_DATA_TEMPR2[19] ), .D(\Z\R_DATA_TEMPR3[19] ), .Y(
        OR4_524_Y));
    OR4 \OR4_R_DATA[28]  (.A(OR4_633_Y), .B(OR4_536_Y), .C(OR4_217_Y), 
        .D(OR4_303_Y), .Y(R_DATA_c[28]));
    OR4 OR4_368 (.A(\Z\R_DATA_TEMPR4[11] ), .B(\Z\R_DATA_TEMPR5[11] ), 
        .C(\Z\R_DATA_TEMPR6[11] ), .D(\Z\R_DATA_TEMPR7[11] ), .Y(
        OR4_368_Y));
    OR4 OR4_712 (.A(OR4_238_Y), .B(OR4_75_Y), .C(OR4_64_Y), .D(
        OR4_514_Y), .Y(OR4_712_Y));
    OR4 OR4_630 (.A(OR4_511_Y), .B(OR4_666_Y), .C(OR4_20_Y), .D(
        OR4_550_Y), .Y(OR4_630_Y));
    OR4 OR4_98 (.A(\Z\R_DATA_TEMPR8[27] ), .B(\Z\R_DATA_TEMPR9[27] ), 
        .C(\Z\R_DATA_TEMPR10[27] ), .D(\Z\R_DATA_TEMPR11[27] ), .Y(
        OR4_98_Y));
    OR4 OR4_321 (.A(\Z\R_DATA_TEMPR0[5] ), .B(\Z\R_DATA_TEMPR1[5] ), 
        .C(\Z\R_DATA_TEMPR2[5] ), .D(\Z\R_DATA_TEMPR3[5] ), .Y(
        OR4_321_Y));
    OR4 OR4_615 (.A(\Z\R_DATA_TEMPR8[75] ), .B(\Z\R_DATA_TEMPR9[75] ), 
        .C(\Z\R_DATA_TEMPR10[75] ), .D(\Z\R_DATA_TEMPR11[75] ), .Y(
        OR4_615_Y));
    OR4 OR4_337 (.A(\Z\R_DATA_TEMPR8[71] ), .B(\Z\R_DATA_TEMPR9[71] ), 
        .C(\Z\R_DATA_TEMPR10[71] ), .D(\Z\R_DATA_TEMPR11[71] ), .Y(
        OR4_337_Y));
    OR4 OR4_130 (.A(\Z\R_DATA_TEMPR16[35] ), .B(\Z\R_DATA_TEMPR17[35] )
        , .C(\Z\R_DATA_TEMPR18[35] ), .D(\Z\R_DATA_TEMPR19[35] ), .Y(
        OR4_130_Y));
    OR2 OR2_25 (.A(\Z\R_DATA_TEMPR20[30] ), .B(\Z\R_DATA_TEMPR21[30] ), 
        .Y(OR2_25_Y));
    OR4 OR4_303 (.A(\Z\R_DATA_TEMPR28[28] ), .B(\Z\R_DATA_TEMPR29[28] )
        , .C(\Z\R_DATA_TEMPR30[28] ), .D(\Z\R_DATA_TEMPR31[28] ), .Y(
        OR4_303_Y));
    OR4 OR4_169 (.A(\Z\R_DATA_TEMPR8[78] ), .B(\Z\R_DATA_TEMPR9[78] ), 
        .C(\Z\R_DATA_TEMPR10[78] ), .D(\Z\R_DATA_TEMPR11[78] ), .Y(
        OR4_169_Y));
    
endmodule


module test2(
       CLK,
       R_ADDR,
       R_EN,
       WBYTE_EN,
       W_ADDR,
       W_DATA,
       W_EN,
       selectt,
       ERRr,
       R_DATA,
       data_64_out,
       error_address,
       error_data,
       error_flag
    );
input  CLK;
input  [13:0] R_ADDR;
input  R_EN;
input  [7:0] WBYTE_EN;
input  [13:0] W_ADDR;
input  [79:0] W_DATA;
input  W_EN;
input  [63:0] selectt;
output ERRr;
output [79:0] R_DATA;
output [63:0] data_64_out;
output [13:0] error_address;
output [63:0] error_data;
output error_flag;

    wire [63:0] data_64_out_net_0;
    wire [7:0] PF_TPSRAM_C0_0_R_DATA;
    wire [7:0] en64_RP2_0_OUTt;
    wire [13:0] R_ADDR_c;
    wire [7:0] WBYTE_EN_c;
    wire [13:0] W_ADDR_c;
    wire [79:0] W_DATA_c;
    wire [63:0] selectt_c;
    wire [79:0] R_DATA_c;
    wire [13:0] error_address_c;
    wire [63:0] error_data_c;
    wire NN_1, GND, VCC, CLK_ibuf_Z, R_EN_c, W_EN_c, ERRr_c, N_24, 
        N_25, N_26, N_27, N_28, N_29, N_30, N_31, N_32, N_33, N_34, 
        N_35, N_36, N_37, N_38, N_39, N_40, N_41, N_42, N_43, N_44, 
        N_45, N_46, N_47, N_48, N_49, N_50, N_51;
    
    OUTBUF \R_DATA_obuf[76]  (.D(R_DATA_c[76]), .PAD(R_DATA[76]));
    OUTBUF \error_data_obuf[2]  (.D(error_data_c[2]), .PAD(
        error_data[2]));
    OUTBUF \data_64_out_obuf[40]  (.D(W_DATA_c[50]), .PAD(
        data_64_out[40]));
    OUTBUF \data_64_out_obuf[36]  (.D(W_DATA_c[44]), .PAD(
        data_64_out[36]));
    INBUF \W_DATA_ibuf[12]  (.PAD(W_DATA[12]), .Y(W_DATA_c[12]));
    INBUF \selectt_ibuf[32]  (.PAD(selectt[32]), .Y(selectt_c[32]));
    INBUF \W_DATA_ibuf[65]  (.PAD(W_DATA[65]), .Y(W_DATA_c[65]));
    INBUF \selectt_ibuf[37]  (.PAD(selectt[37]), .Y(selectt_c[37]));
    OUTBUF \error_data_obuf[18]  (.D(error_data_c[18]), .PAD(
        error_data[18]));
    OUTBUF \error_address_obuf[0]  (.D(error_address_c[0]), .PAD(
        error_address[0]));
    INBUF \selectt_ibuf[41]  (.PAD(selectt[41]), .Y(selectt_c[41]));
    INBUF \selectt_ibuf[36]  (.PAD(selectt[36]), .Y(selectt_c[36]));
    OUTBUF \data_64_out_obuf[51]  (.D(W_DATA_c[63]), .PAD(
        data_64_out[51]));
    test6_for_compare test6_for_compare_0 (.error_data_c({
        error_data_c[63], error_data_c[62], error_data_c[61], 
        error_data_c[60], error_data_c[59], error_data_c[58], 
        error_data_c[57], error_data_c[56], error_data_c[55], 
        error_data_c[54], error_data_c[53], error_data_c[52], 
        error_data_c[51], error_data_c[50], error_data_c[49], 
        error_data_c[48], error_data_c[47], error_data_c[46], 
        error_data_c[45], error_data_c[44], error_data_c[43], 
        error_data_c[42], error_data_c[41], error_data_c[40], 
        error_data_c[39], error_data_c[38], error_data_c[37], 
        error_data_c[36], error_data_c[35], error_data_c[34], 
        error_data_c[33], error_data_c[32], error_data_c[31], 
        error_data_c[30], error_data_c[29], error_data_c[28], 
        error_data_c[27], error_data_c[26], error_data_c[25], 
        error_data_c[24], error_data_c[23], error_data_c[22], 
        error_data_c[21], error_data_c[20], error_data_c[19], 
        error_data_c[18], error_data_c[17], error_data_c[16], 
        error_data_c[15], error_data_c[14], error_data_c[13], 
        error_data_c[12], error_data_c[11], error_data_c[10], 
        error_data_c[9], error_data_c[8], error_data_c[7], 
        error_data_c[6], error_data_c[5], error_data_c[4], 
        error_data_c[3], error_data_c[2], error_data_c[1], 
        error_data_c[0]}), .data_64_out_net_0({data_64_out_net_0[63], 
        data_64_out_net_0[62], data_64_out_net_0[61], 
        data_64_out_net_0[60], data_64_out_net_0[59], 
        data_64_out_net_0[58], data_64_out_net_0[57], 
        data_64_out_net_0[56], data_64_out_net_0[55], 
        data_64_out_net_0[54], data_64_out_net_0[53], 
        data_64_out_net_0[52], data_64_out_net_0[51], 
        data_64_out_net_0[50], data_64_out_net_0[49], 
        data_64_out_net_0[48], data_64_out_net_0[47], 
        data_64_out_net_0[46], data_64_out_net_0[45], 
        data_64_out_net_0[44], data_64_out_net_0[43], 
        data_64_out_net_0[42], data_64_out_net_0[41], 
        data_64_out_net_0[40], data_64_out_net_0[39], 
        data_64_out_net_0[38], data_64_out_net_0[37], 
        data_64_out_net_0[36], data_64_out_net_0[35], 
        data_64_out_net_0[34], data_64_out_net_0[33], 
        data_64_out_net_0[32], data_64_out_net_0[31], 
        data_64_out_net_0[30], data_64_out_net_0[29], 
        data_64_out_net_0[28], data_64_out_net_0[27], 
        data_64_out_net_0[26], data_64_out_net_0[25], 
        data_64_out_net_0[24], data_64_out_net_0[23], 
        data_64_out_net_0[22], data_64_out_net_0[21], 
        data_64_out_net_0[20], data_64_out_net_0[19], 
        data_64_out_net_0[18], data_64_out_net_0[17], 
        data_64_out_net_0[16], data_64_out_net_0[15], 
        data_64_out_net_0[14], data_64_out_net_0[13], 
        data_64_out_net_0[12], data_64_out_net_0[11], 
        data_64_out_net_0[10], data_64_out_net_0[9], 
        data_64_out_net_0[8], data_64_out_net_0[7], 
        data_64_out_net_0[6], data_64_out_net_0[5], 
        data_64_out_net_0[4], data_64_out_net_0[3], 
        data_64_out_net_0[2], data_64_out_net_0[1], 
        data_64_out_net_0[0]}), .error_address_c({error_address_c[13], 
        error_address_c[12], error_address_c[11], error_address_c[10], 
        error_address_c[9], error_address_c[8], error_address_c[7], 
        error_address_c[6], error_address_c[5], error_address_c[4], 
        error_address_c[3], error_address_c[2], error_address_c[1], 
        error_address_c[0]}), .R_ADDR_c({R_ADDR_c[13], R_ADDR_c[12], 
        R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0]}), .ERRr_c(
        ERRr_c));
    OUTBUF \error_data_obuf[45]  (.D(error_data_c[45]), .PAD(
        error_data[45]));
    INBUF \W_DATA_ibuf[60]  (.PAD(W_DATA[60]), .Y(W_DATA_c[60]));
    OUTBUF \error_data_obuf[36]  (.D(error_data_c[36]), .PAD(
        error_data[36]));
    OUTBUF \error_data_obuf[1]  (.D(error_data_c[1]), .PAD(
        error_data[1]));
    INBUF \W_DATA_ibuf[32]  (.PAD(W_DATA[32]), .Y(W_DATA_c[32]));
    OUTBUF \data_64_out_obuf[37]  (.D(W_DATA_c[45]), .PAD(
        data_64_out[37]));
    OUTBUF \data_64_out_obuf[24]  (.D(W_DATA_c[30]), .PAD(
        data_64_out[24]));
    INBUF \selectt_ibuf[18]  (.PAD(selectt[18]), .Y(selectt_c[18]));
    OUTBUF \error_data_obuf[32]  (.D(error_data_c[32]), .PAD(
        error_data[32]));
    INBUF \selectt_ibuf[55]  (.PAD(selectt[55]), .Y(selectt_c[55]));
    INBUF \selectt_ibuf[10]  (.PAD(selectt[10]), .Y(selectt_c[10]));
    INBUF \selectt_ibuf[0]  (.PAD(selectt[0]), .Y(selectt_c[0]));
    OUTBUF \error_data_obuf[44]  (.D(error_data_c[44]), .PAD(
        error_data[44]));
    INBUF \W_DATA_ibuf[18]  (.PAD(W_DATA[18]), .Y(W_DATA_c[18]));
    OUTBUF \error_data_obuf[20]  (.D(error_data_c[20]), .PAD(
        error_data[20]));
    INBUF \W_ADDR_ibuf[5]  (.PAD(W_ADDR[5]), .Y(W_ADDR_c[5]));
    OUTBUF \R_DATA_obuf[45]  (.D(R_DATA_c[45]), .PAD(R_DATA[45]));
    OUTBUF \data_64_out_obuf[11]  (.D(W_DATA_c[13]), .PAD(
        data_64_out[11]));
    INBUF \W_DATA_ibuf[16]  (.PAD(W_DATA[16]), .Y(W_DATA_c[16]));
    INBUF \W_ADDR_ibuf[12]  (.PAD(W_ADDR[12]), .Y(W_ADDR_c[12]));
    INBUF \W_DATA_ibuf[45]  (.PAD(W_DATA[45]), .Y(W_DATA_c[45]));
    OUTBUF \data_64_out_obuf[4]  (.D(W_DATA_c[4]), .PAD(data_64_out[4])
        );
    INBUF \W_DATA_ibuf[38]  (.PAD(W_DATA[38]), .Y(W_DATA_c[38]));
    INBUF \W_DATA_ibuf[21]  (.PAD(W_DATA[21]), .Y(W_DATA_c[21]));
    OUTBUF \R_DATA_obuf[37]  (.D(R_DATA_c[37]), .PAD(R_DATA[37]));
    INBUF \W_DATA_ibuf[51]  (.PAD(W_DATA[51]), .Y(W_DATA_c[51]));
    INBUF \W_DATA_ibuf[73]  (.PAD(W_DATA[73]), .Y(W_DATA_c[73]));
    OUTBUF \data_64_out_obuf[41]  (.D(W_DATA_c[51]), .PAD(
        data_64_out[41]));
    INBUF \W_DATA_ibuf[40]  (.PAD(W_DATA[40]), .Y(W_DATA_c[40]));
    INBUF \W_DATA_ibuf[36]  (.PAD(W_DATA[36]), .Y(W_DATA_c[36]));
    INBUF \WBYTE_EN_ibuf[5]  (.PAD(WBYTE_EN[5]), .Y(WBYTE_EN_c[5]));
    INBUF \selectt_ibuf[14]  (.PAD(selectt[14]), .Y(selectt_c[14]));
    OUTBUF \R_DATA_obuf[43]  (.D(R_DATA_c[43]), .PAD(R_DATA[43]));
    INBUF \W_ADDR_ibuf[3]  (.PAD(W_ADDR[3]), .Y(W_ADDR_c[3]));
    INBUF \W_ADDR_ibuf[2]  (.PAD(W_ADDR[2]), .Y(W_ADDR_c[2]));
    OUTBUF \error_address_obuf[9]  (.D(error_address_c[9]), .PAD(
        error_address[9]));
    OUTBUF \R_DATA_obuf[30]  (.D(R_DATA_c[30]), .PAD(R_DATA[30]));
    OUTBUF \data_64_out_obuf[5]  (.D(W_DATA_c[5]), .PAD(data_64_out[5])
        );
    OUTBUF \error_data_obuf[23]  (.D(error_data_c[23]), .PAD(
        error_data[23]));
    en64_RP2 en64_RP2_0 (.en64_RP2_0_OUTt({en64_RP2_0_OUTt[7], 
        en64_RP2_0_OUTt[6], en64_RP2_0_OUTt[5], en64_RP2_0_OUTt[4], 
        en64_RP2_0_OUTt[3], en64_RP2_0_OUTt[2], en64_RP2_0_OUTt[1], 
        en64_RP2_0_OUTt[0]}), .W_DATA_c({W_DATA_c[77], W_DATA_c[76], 
        W_DATA_c[75], W_DATA_c[74], W_DATA_c[73], W_DATA_c[72], 
        W_DATA_c[71], W_DATA_c[70], N_37, N_36, W_DATA_c[67], 
        W_DATA_c[66], W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], 
        W_DATA_c[62], W_DATA_c[61], W_DATA_c[60], N_35, N_34, 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], N_33, 
        N_32, W_DATA_c[47], W_DATA_c[46], W_DATA_c[45], W_DATA_c[44], 
        W_DATA_c[43], W_DATA_c[42], W_DATA_c[41], W_DATA_c[40], N_31, 
        N_30, W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], N_29, 
        N_28, W_DATA_c[27], W_DATA_c[26], W_DATA_c[25], W_DATA_c[24], 
        W_DATA_c[23], W_DATA_c[22], W_DATA_c[21], W_DATA_c[20], N_27, 
        N_26, W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], N_25, 
        N_24, W_DATA_c[7], W_DATA_c[6], W_DATA_c[5], W_DATA_c[4], 
        W_DATA_c[3], W_DATA_c[2], W_DATA_c[1], W_DATA_c[0]}));
    INBUF \selectt_ibuf[4]  (.PAD(selectt[4]), .Y(selectt_c[4]));
    OUTBUF \error_address_obuf[7]  (.D(error_address_c[7]), .PAD(
        error_address[7]));
    OUTBUF \R_DATA_obuf[59]  (.D(R_DATA_c[59]), .PAD(R_DATA[59]));
    OUTBUF \data_64_out_obuf[6]  (.D(W_DATA_c[6]), .PAD(data_64_out[6])
        );
    OUTBUF \error_data_obuf[58]  (.D(error_data_c[58]), .PAD(
        error_data[58]));
    OUTBUF \R_DATA_obuf[2]  (.D(R_DATA_c[2]), .PAD(R_DATA[2]));
    OUTBUF \R_DATA_obuf[44]  (.D(R_DATA_c[44]), .PAD(R_DATA[44]));
    OUTBUF \data_64_out_obuf[58]  (.D(W_DATA_c[72]), .PAD(
        data_64_out[58]));
    OUTBUF \R_DATA_obuf[56]  (.D(R_DATA_c[56]), .PAD(R_DATA[56]));
    OUTBUF \R_DATA_obuf[15]  (.D(R_DATA_c[15]), .PAD(R_DATA[15]));
    INBUF \R_ADDR_ibuf[6]  (.PAD(R_ADDR[6]), .Y(R_ADDR_c[6]));
    OUTBUF \R_DATA_obuf[25]  (.D(R_DATA_c[25]), .PAD(R_DATA[25]));
    OUTBUF \error_data_obuf[3]  (.D(error_data_c[3]), .PAD(
        error_data[3]));
    OUTBUF \error_data_obuf[7]  (.D(error_data_c[7]), .PAD(
        error_data[7]));
    OUTBUF \R_DATA_obuf[67]  (.D(R_DATA_c[67]), .PAD(R_DATA[67]));
    INBUF \selectt_ibuf[62]  (.PAD(selectt[62]), .Y(selectt_c[62]));
    OUTBUF \error_data_obuf[41]  (.D(error_data_c[41]), .PAD(
        error_data[41]));
    INBUF \W_DATA_ibuf[11]  (.PAD(W_DATA[11]), .Y(W_DATA_c[11]));
    OUTBUF \error_data_obuf[29]  (.D(error_data_c[29]), .PAD(
        error_data[29]));
    INBUF W_EN_ibuf (.PAD(W_EN), .Y(W_EN_c));
    INBUF \selectt_ibuf[39]  (.PAD(selectt[39]), .Y(selectt_c[39]));
    OUTBUF \R_DATA_obuf[13]  (.D(R_DATA_c[13]), .PAD(R_DATA[13]));
    OUTBUF \data_64_out_obuf[33]  (.D(W_DATA_c[41]), .PAD(
        data_64_out[33]));
    OUTBUF \R_DATA_obuf[60]  (.D(R_DATA_c[60]), .PAD(R_DATA[60]));
    OUTBUF \R_DATA_obuf[23]  (.D(R_DATA_c[23]), .PAD(R_DATA[23]));
    OUTBUF \R_DATA_obuf[32]  (.D(R_DATA_c[32]), .PAD(R_DATA[32]));
    de_v1 de_v1_0 (.data_64_out_net_0({data_64_out_net_0[63], 
        data_64_out_net_0[62], data_64_out_net_0[61], 
        data_64_out_net_0[60], data_64_out_net_0[59], 
        data_64_out_net_0[58], data_64_out_net_0[57], 
        data_64_out_net_0[56], data_64_out_net_0[55], 
        data_64_out_net_0[54], data_64_out_net_0[53], 
        data_64_out_net_0[52], data_64_out_net_0[51], 
        data_64_out_net_0[50], data_64_out_net_0[49], 
        data_64_out_net_0[48], data_64_out_net_0[47], 
        data_64_out_net_0[46], data_64_out_net_0[45], 
        data_64_out_net_0[44], data_64_out_net_0[43], 
        data_64_out_net_0[42], data_64_out_net_0[41], 
        data_64_out_net_0[40], data_64_out_net_0[39], 
        data_64_out_net_0[38], data_64_out_net_0[37], 
        data_64_out_net_0[36], data_64_out_net_0[35], 
        data_64_out_net_0[34], data_64_out_net_0[33], 
        data_64_out_net_0[32], data_64_out_net_0[31], 
        data_64_out_net_0[30], data_64_out_net_0[29], 
        data_64_out_net_0[28], data_64_out_net_0[27], 
        data_64_out_net_0[26], data_64_out_net_0[25], 
        data_64_out_net_0[24], data_64_out_net_0[23], 
        data_64_out_net_0[22], data_64_out_net_0[21], 
        data_64_out_net_0[20], data_64_out_net_0[19], 
        data_64_out_net_0[18], data_64_out_net_0[17], 
        data_64_out_net_0[16], data_64_out_net_0[15], 
        data_64_out_net_0[14], data_64_out_net_0[13], 
        data_64_out_net_0[12], data_64_out_net_0[11], 
        data_64_out_net_0[10], data_64_out_net_0[9], 
        data_64_out_net_0[8], data_64_out_net_0[7], 
        data_64_out_net_0[6], data_64_out_net_0[5], 
        data_64_out_net_0[4], data_64_out_net_0[3], 
        data_64_out_net_0[2], data_64_out_net_0[1], 
        data_64_out_net_0[0]}), .PF_TPSRAM_C0_0_R_DATA({
        PF_TPSRAM_C0_0_R_DATA[7], PF_TPSRAM_C0_0_R_DATA[6], 
        PF_TPSRAM_C0_0_R_DATA[5], PF_TPSRAM_C0_0_R_DATA[4], 
        PF_TPSRAM_C0_0_R_DATA[3], PF_TPSRAM_C0_0_R_DATA[2], 
        PF_TPSRAM_C0_0_R_DATA[1], PF_TPSRAM_C0_0_R_DATA[0]}), .ERRr_c(
        ERRr_c));
    OUTBUF \data_64_out_obuf[18]  (.D(W_DATA_c[22]), .PAD(
        data_64_out[18]));
    OUTBUF \R_DATA_obuf[48]  (.D(R_DATA_c[48]), .PAD(R_DATA[48]));
    INBUF \WBYTE_EN_ibuf[7]  (.PAD(WBYTE_EN[7]), .Y(WBYTE_EN_c[7]));
    OUTBUF \error_data_obuf[17]  (.D(error_data_c[17]), .PAD(
        error_data[17]));
    OUTBUF \error_address_obuf[8]  (.D(error_address_c[8]), .PAD(
        error_address[8]));
    INBUF \W_DATA_ibuf[31]  (.PAD(W_DATA[31]), .Y(W_DATA_c[31]));
    INBUF \W_DATA_ibuf[23]  (.PAD(W_DATA[23]), .Y(W_DATA_c[23]));
    OUTBUF \data_64_out_obuf[20]  (.D(W_DATA_c[24]), .PAD(
        data_64_out[20]));
    OUTBUF \R_DATA_obuf[4]  (.D(R_DATA_c[4]), .PAD(R_DATA[4]));
    INBUF \R_ADDR_ibuf[9]  (.PAD(R_ADDR[9]), .Y(R_ADDR_c[9]));
    INBUF \W_DATA_ibuf[53]  (.PAD(W_DATA[53]), .Y(W_DATA_c[53]));
    INBUF \W_DATA_ibuf[1]  (.PAD(W_DATA[1]), .Y(W_DATA_c[1]));
    OUTBUF \R_DATA_obuf[6]  (.D(R_DATA_c[6]), .PAD(R_DATA[6]));
    INBUF \selectt_ibuf[52]  (.PAD(selectt[52]), .Y(selectt_c[52]));
    INBUF \selectt_ibuf[43]  (.PAD(selectt[43]), .Y(selectt_c[43]));
    INBUF \selectt_ibuf[57]  (.PAD(selectt[57]), .Y(selectt_c[57]));
    INBUF \selectt_ibuf[56]  (.PAD(selectt[56]), .Y(selectt_c[56]));
    OUTBUF \data_64_out_obuf[48]  (.D(W_DATA_c[60]), .PAD(
        data_64_out[48]));
    OUTBUF \R_DATA_obuf[41]  (.D(R_DATA_c[41]), .PAD(R_DATA[41]));
    INBUF \R_ADDR_ibuf[10]  (.PAD(R_ADDR[10]), .Y(R_ADDR_c[10]));
    OUTBUF \R_DATA_obuf[14]  (.D(R_DATA_c[14]), .PAD(R_DATA[14]));
    OUTBUF \R_DATA_obuf[24]  (.D(R_DATA_c[24]), .PAD(R_DATA[24]));
    INBUF \selectt_ibuf[38]  (.PAD(selectt[38]), .Y(selectt_c[38]));
    INBUF \selectt_ibuf[30]  (.PAD(selectt[30]), .Y(selectt_c[30]));
    INBUF \selectt_ibuf[1]  (.PAD(selectt[1]), .Y(selectt_c[1]));
    INBUF \W_ADDR_ibuf[7]  (.PAD(W_ADDR[7]), .Y(W_ADDR_c[7]));
    OUTBUF \data_64_out_obuf[3]  (.D(W_DATA_c[3]), .PAD(data_64_out[3])
        );
    INBUF \selectt_ibuf[11]  (.PAD(selectt[11]), .Y(selectt_c[11]));
    OUTBUF \R_DATA_obuf[62]  (.D(R_DATA_c[62]), .PAD(R_DATA[62]));
    OUTBUF \R_DATA_obuf[18]  (.D(R_DATA_c[18]), .PAD(R_DATA[18]));
    INBUF \W_DATA_ibuf[74]  (.PAD(W_DATA[74]), .Y(W_DATA_c[74]));
    OUTBUF \R_DATA_obuf[28]  (.D(R_DATA_c[28]), .PAD(R_DATA[28]));
    OUTBUF \error_data_obuf[46]  (.D(error_data_c[46]), .PAD(
        error_data[46]));
    INBUF \W_ADDR_ibuf[8]  (.PAD(W_ADDR[8]), .Y(W_ADDR_c[8]));
    INBUF \selectt_ibuf[34]  (.PAD(selectt[34]), .Y(selectt_c[34]));
    OUTBUF \data_64_out_obuf[21]  (.D(W_DATA_c[25]), .PAD(
        data_64_out[21]));
    INBUF \W_DATA_ibuf[13]  (.PAD(W_DATA[13]), .Y(W_DATA_c[13]));
    OUTBUF \data_64_out_obuf[60]  (.D(W_DATA_c[74]), .PAD(
        data_64_out[60]));
    OUTBUF \error_data_obuf[42]  (.D(error_data_c[42]), .PAD(
        error_data[42]));
    OUTBUF \data_64_out_obuf[0]  (.D(W_DATA_c[0]), .PAD(data_64_out[0])
        );
    OUTBUF \data_64_out_obuf[39]  (.D(W_DATA_c[47]), .PAD(
        data_64_out[39]));
    OUTBUF \R_DATA_obuf[11]  (.D(R_DATA_c[11]), .PAD(R_DATA[11]));
    INBUF \R_ADDR_ibuf[13]  (.PAD(R_ADDR[13]), .Y(R_ADDR_c[13]));
    OUTBUF \R_DATA_obuf[21]  (.D(R_DATA_c[21]), .PAD(R_DATA[21]));
    INBUF \W_DATA_ibuf[33]  (.PAD(W_DATA[33]), .Y(W_DATA_c[33]));
    OUTBUF \error_data_obuf[57]  (.D(error_data_c[57]), .PAD(
        error_data[57]));
    OUTBUF \data_64_out_obuf[55]  (.D(W_DATA_c[67]), .PAD(
        data_64_out[55]));
    OUTBUF \error_data_obuf[10]  (.D(error_data_c[10]), .PAD(
        error_data[10]));
    OUTBUF \data_64_out_obuf[56]  (.D(W_DATA_c[70]), .PAD(
        data_64_out[56]));
    OUTBUF \data_64_out_obuf[1]  (.D(W_DATA_c[1]), .PAD(data_64_out[1])
        );
    OUTBUF \error_address_obuf[6]  (.D(error_address_c[6]), .PAD(
        error_address[6]));
    OUTBUF \error_address_obuf[11]  (.D(error_address_c[11]), .PAD(
        error_address[11]));
    INBUF \selectt_ibuf[25]  (.PAD(selectt[25]), .Y(selectt_c[25]));
    INBUF \W_DATA_ibuf[69]  (.PAD(W_DATA[69]), .Y(W_DATA_c[69]));
    OUTBUF \error_data_obuf[25]  (.D(error_data_c[25]), .PAD(
        error_data[25]));
    OUTBUF ERRr_obuf (.D(ERRr_c), .PAD(ERRr));
    OUTBUF \data_64_out_obuf[57]  (.D(W_DATA_c[71]), .PAD(
        data_64_out[57]));
    OUTBUF \data_64_out_obuf[15]  (.D(W_DATA_c[17]), .PAD(
        data_64_out[15]));
    OUTBUF \error_data_obuf[24]  (.D(error_data_c[24]), .PAD(
        error_data[24]));
    OUTBUF \R_DATA_obuf[35]  (.D(R_DATA_c[35]), .PAD(R_DATA[35]));
    OUTBUF \data_64_out_obuf[2]  (.D(W_DATA_c[2]), .PAD(data_64_out[2])
        );
    INBUF \W_DATA_ibuf[6]  (.PAD(W_DATA[6]), .Y(W_DATA_c[6]));
    INBUF \selectt_ibuf[59]  (.PAD(selectt[59]), .Y(selectt_c[59]));
    OUTBUF \data_64_out_obuf[61]  (.D(W_DATA_c[75]), .PAD(
        data_64_out[61]));
    OUTBUF \data_64_out_obuf[16]  (.D(W_DATA_c[20]), .PAD(
        data_64_out[16]));
    OUTBUF \error_data_obuf[38]  (.D(error_data_c[38]), .PAD(
        error_data[38]));
    OUTBUF \error_data_obuf[13]  (.D(error_data_c[13]), .PAD(
        error_data[13]));
    INBUF \W_DATA_ibuf[24]  (.PAD(W_DATA[24]), .Y(W_DATA_c[24]));
    INBUF \selectt_ibuf[60]  (.PAD(selectt[60]), .Y(selectt_c[60]));
    OUTBUF \data_64_out_obuf[45]  (.D(W_DATA_c[55]), .PAD(
        data_64_out[45]));
    OUTBUF \R_DATA_obuf[49]  (.D(R_DATA_c[49]), .PAD(R_DATA[49]));
    INBUF \W_DATA_ibuf[54]  (.PAD(W_DATA[54]), .Y(W_DATA_c[54]));
    INBUF \W_DATA_ibuf[67]  (.PAD(W_DATA[67]), .Y(W_DATA_c[67]));
    INBUF \W_ADDR_ibuf[6]  (.PAD(W_ADDR[6]), .Y(W_ADDR_c[6]));
    OUTBUF \R_DATA_obuf[33]  (.D(R_DATA_c[33]), .PAD(R_DATA[33]));
    OUTBUF \data_64_out_obuf[46]  (.D(W_DATA_c[56]), .PAD(
        data_64_out[46]));
    INBUF \W_DATA_ibuf[4]  (.PAD(W_DATA[4]), .Y(W_DATA_c[4]));
    OUTBUF \data_64_out_obuf[17]  (.D(W_DATA_c[21]), .PAD(
        data_64_out[17]));
    INBUF \W_DATA_ibuf[49]  (.PAD(W_DATA[49]), .Y(W_DATA_c[49]));
    INBUF \selectt_ibuf[3]  (.PAD(selectt[3]), .Y(selectt_c[3]));
    OUTBUF \data_64_out_obuf[28]  (.D(W_DATA_c[34]), .PAD(
        data_64_out[28]));
    OUTBUF \R_DATA_obuf[46]  (.D(R_DATA_c[46]), .PAD(R_DATA[46]));
    OUTBUF \error_data_obuf[60]  (.D(error_data_c[60]), .PAD(
        error_data[60]));
    OUTBUF \data_64_out_obuf[8]  (.D(W_DATA_c[10]), .PAD(
        data_64_out[8]));
    INBUF \W_DATA_ibuf[75]  (.PAD(W_DATA[75]), .Y(W_DATA_c[75]));
    INBUF \R_ADDR_ibuf[7]  (.PAD(R_ADDR[7]), .Y(R_ADDR_c[7]));
    INBUF \selectt_ibuf[58]  (.PAD(selectt[58]), .Y(selectt_c[58]));
    OUTBUF \error_address_obuf[4]  (.D(error_address_c[4]), .PAD(
        error_address[4]));
    INBUF \selectt_ibuf[50]  (.PAD(selectt[50]), .Y(selectt_c[50]));
    OUTBUF \data_64_out_obuf[47]  (.D(W_DATA_c[57]), .PAD(
        data_64_out[47]));
    INBUF \W_DATA_ibuf[2]  (.PAD(W_DATA[2]), .Y(W_DATA_c[2]));
    OUTBUF \error_address_obuf[1]  (.D(error_address_c[1]), .PAD(
        error_address[1]));
    OUTBUF \data_64_out_obuf[32]  (.D(W_DATA_c[40]), .PAD(
        data_64_out[32]));
    INBUF \W_DATA_ibuf[70]  (.PAD(W_DATA[70]), .Y(W_DATA_c[70]));
    OUTBUF \error_data_obuf[19]  (.D(error_data_c[19]), .PAD(
        error_data[19]));
    OUTBUF \R_DATA_obuf[65]  (.D(R_DATA_c[65]), .PAD(R_DATA[65]));
    OUTBUF \R_DATA_obuf[34]  (.D(R_DATA_c[34]), .PAD(R_DATA[34]));
    INBUF \selectt_ibuf[31]  (.PAD(selectt[31]), .Y(selectt_c[31]));
    OUTBUF \error_data_obuf[50]  (.D(error_data_c[50]), .PAD(
        error_data[50]));
    INBUF \selectt_ibuf[13]  (.PAD(selectt[13]), .Y(selectt_c[13]));
    INBUF \W_DATA_ibuf[47]  (.PAD(W_DATA[47]), .Y(W_DATA_c[47]));
    OUTBUF \error_address_obuf[2]  (.D(error_address_c[2]), .PAD(
        error_address[2]));
    OUTBUF \error_data_obuf[63]  (.D(error_data_c[63]), .PAD(
        error_data[63]));
    INBUF \W_DATA_ibuf[14]  (.PAD(W_DATA[14]), .Y(W_DATA_c[14]));
    OUTBUF \R_DATA_obuf[63]  (.D(R_DATA_c[63]), .PAD(R_DATA[63]));
    OUTBUF \R_DATA_obuf[19]  (.D(R_DATA_c[19]), .PAD(R_DATA[19]));
    INBUF \selectt_ibuf[54]  (.PAD(selectt[54]), .Y(selectt_c[54]));
    OUTBUF \R_DATA_obuf[29]  (.D(R_DATA_c[29]), .PAD(R_DATA[29]));
    INBUF \R_ADDR_ibuf[4]  (.PAD(R_ADDR[4]), .Y(R_ADDR_c[4]));
    OUTBUF \error_data_obuf[21]  (.D(error_data_c[21]), .PAD(
        error_data[21]));
    OUTBUF \error_address_obuf[10]  (.D(error_address_c[10]), .PAD(
        error_address[10]));
    INBUF \selectt_ibuf[2]  (.PAD(selectt[2]), .Y(selectt_c[2]));
    OUTBUF \R_DATA_obuf[38]  (.D(R_DATA_c[38]), .PAD(R_DATA[38]));
    OUTBUF \R_DATA_obuf[16]  (.D(R_DATA_c[16]), .PAD(R_DATA[16]));
    INBUF \W_DATA_ibuf[34]  (.PAD(W_DATA[34]), .Y(W_DATA_c[34]));
    INBUF \selectt_ibuf[22]  (.PAD(selectt[22]), .Y(selectt_c[22]));
    OUTBUF \R_DATA_obuf[26]  (.D(R_DATA_c[26]), .PAD(R_DATA[26]));
    OUTBUF \error_data_obuf[53]  (.D(error_data_c[53]), .PAD(
        error_data[53]));
    INBUF \selectt_ibuf[27]  (.PAD(selectt[27]), .Y(selectt_c[27]));
    OUTBUF \data_64_out_obuf[53]  (.D(W_DATA_c[65]), .PAD(
        data_64_out[53]));
    INBUF \selectt_ibuf[26]  (.PAD(selectt[26]), .Y(selectt_c[26]));
    GND GND_Z (.Y(GND));
    OUTBUF \R_DATA_obuf[64]  (.D(R_DATA_c[64]), .PAD(R_DATA[64]));
    OUTBUF \R_DATA_obuf[31]  (.D(R_DATA_c[31]), .PAD(R_DATA[31]));
    INBUF \W_DATA_ibuf[7]  (.PAD(W_DATA[7]), .Y(W_DATA_c[7]));
    INBUF \W_DATA_ibuf[25]  (.PAD(W_DATA[25]), .Y(W_DATA_c[25]));
    VCC VCC_Z (.Y(VCC));
    INBUF \W_DATA_ibuf[55]  (.PAD(W_DATA[55]), .Y(W_DATA_c[55]));
    INBUF \W_DATA_ibuf[20]  (.PAD(W_DATA[20]), .Y(W_DATA_c[20]));
    OUTBUF \data_64_out_obuf[13]  (.D(W_DATA_c[15]), .PAD(
        data_64_out[13]));
    INBUF CLK_ibuf (.PAD(CLK), .Y(CLK_ibuf_Z));
    INBUF \W_DATA_ibuf[50]  (.PAD(W_DATA[50]), .Y(W_DATA_c[50]));
    OUTBUF \R_DATA_obuf[77]  (.D(R_DATA_c[77]), .PAD(R_DATA[77]));
    OUTBUF \error_data_obuf[37]  (.D(error_data_c[37]), .PAD(
        error_data[37]));
    OUTBUF \error_data_obuf[59]  (.D(error_data_c[59]), .PAD(
        error_data[59]));
    OUTBUF \R_DATA_obuf[68]  (.D(R_DATA_c[68]), .PAD(R_DATA[68]));
    OUTBUF \data_64_out_obuf[43]  (.D(W_DATA_c[53]), .PAD(
        data_64_out[43]));
    OUTBUF \R_DATA_obuf[70]  (.D(R_DATA_c[70]), .PAD(R_DATA[70]));
    OUTBUF \data_64_out_obuf[25]  (.D(W_DATA_c[31]), .PAD(
        data_64_out[25]));
    INBUF \WBYTE_EN_ibuf[4]  (.PAD(WBYTE_EN[4]), .Y(WBYTE_EN_c[4]));
    OUTBUF \error_data_obuf[6]  (.D(error_data_c[6]), .PAD(
        error_data[6]));
    OUTBUF \error_data_obuf[26]  (.D(error_data_c[26]), .PAD(
        error_data[26]));
    OUTBUF \data_64_out_obuf[26]  (.D(W_DATA_c[32]), .PAD(
        data_64_out[26]));
    INBUF \W_DATA_ibuf[62]  (.PAD(W_DATA[62]), .Y(W_DATA_c[62]));
    INBUF \selectt_ibuf[61]  (.PAD(selectt[61]), .Y(selectt_c[61]));
    OUTBUF \R_DATA_obuf[61]  (.D(R_DATA_c[61]), .PAD(R_DATA[61]));
    INBUF \selectt_ibuf[6]  (.PAD(selectt[6]), .Y(selectt_c[6]));
    OUTBUF \error_data_obuf[22]  (.D(error_data_c[22]), .PAD(
        error_data[22]));
    OUTBUF \error_data_obuf[15]  (.D(error_data_c[15]), .PAD(
        error_data[15]));
    INBUF \selectt_ibuf[45]  (.PAD(selectt[45]), .Y(selectt_c[45]));
    PF_TPSRAM_C0 PF_TPSRAM_C0_0 (.R_ADDR_c({R_ADDR_c[13], R_ADDR_c[12], 
        R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0]}), 
        .W_ADDR_c({W_ADDR_c[13], W_ADDR_c[12], W_ADDR_c[11], 
        W_ADDR_c[10], W_ADDR_c[9], W_ADDR_c[8], W_ADDR_c[7], 
        W_ADDR_c[6], W_ADDR_c[5], W_ADDR_c[4], W_ADDR_c[3], 
        W_ADDR_c[2], W_ADDR_c[1], W_ADDR_c[0]}), 
        .PF_TPSRAM_C0_0_R_DATA({PF_TPSRAM_C0_0_R_DATA[7], 
        PF_TPSRAM_C0_0_R_DATA[6], PF_TPSRAM_C0_0_R_DATA[5], 
        PF_TPSRAM_C0_0_R_DATA[4], PF_TPSRAM_C0_0_R_DATA[3], 
        PF_TPSRAM_C0_0_R_DATA[2], PF_TPSRAM_C0_0_R_DATA[1], 
        PF_TPSRAM_C0_0_R_DATA[0]}), .en64_RP2_0_OUTt({
        en64_RP2_0_OUTt[7], en64_RP2_0_OUTt[6], en64_RP2_0_OUTt[5], 
        en64_RP2_0_OUTt[4], en64_RP2_0_OUTt[3], en64_RP2_0_OUTt[2], 
        en64_RP2_0_OUTt[1], en64_RP2_0_OUTt[0]}), .CLK(NN_1), .R_EN_c(
        R_EN_c), .W_EN_c(W_EN_c));
    OUTBUF \data_64_out_obuf[59]  (.D(W_DATA_c[73]), .PAD(
        data_64_out[59]));
    INBUF \W_ADDR_ibuf[10]  (.PAD(W_ADDR[10]), .Y(W_ADDR_c[10]));
    INBUF \WBYTE_EN_ibuf[3]  (.PAD(WBYTE_EN[3]), .Y(WBYTE_EN_c[3]));
    INBUF \W_DATA_ibuf[15]  (.PAD(W_DATA[15]), .Y(W_DATA_c[15]));
    OUTBUF \error_data_obuf[48]  (.D(error_data_c[48]), .PAD(
        error_data[48]));
    OUTBUF \data_64_out_obuf[27]  (.D(W_DATA_c[33]), .PAD(
        data_64_out[27]));
    OUTBUF \error_data_obuf[14]  (.D(error_data_c[14]), .PAD(
        error_data[14]));
    INBUF \W_DATA_ibuf[10]  (.PAD(W_DATA[10]), .Y(W_DATA_c[10]));
    INBUF \selectt_ibuf[33]  (.PAD(selectt[33]), .Y(selectt_c[33]));
    INBUF \W_DATA_ibuf[68]  (.PAD(W_DATA[68]), .Y(W_DATA_c[68]));
    INBUF \selectt_ibuf[51]  (.PAD(selectt[51]), .Y(selectt_c[51]));
    OUTBUF \data_64_out_obuf[7]  (.D(W_DATA_c[7]), .PAD(data_64_out[7])
        );
    OUTBUF \data_64_out_obuf[34]  (.D(W_DATA_c[42]), .PAD(
        data_64_out[34]));
    INBUF \W_DATA_ibuf[35]  (.PAD(W_DATA[35]), .Y(W_DATA_c[35]));
    INBUF \R_ADDR_ibuf[11]  (.PAD(R_ADDR[11]), .Y(R_ADDR_c[11]));
    INBUF \WBYTE_EN_ibuf[6]  (.PAD(WBYTE_EN[6]), .Y(WBYTE_EN_c[6]));
    INBUF \W_DATA_ibuf[66]  (.PAD(W_DATA[66]), .Y(W_DATA_c[66]));
    INBUF \selectt_ibuf[5]  (.PAD(selectt[5]), .Y(selectt_c[5]));
    OUTBUF \R_DATA_obuf[72]  (.D(R_DATA_c[72]), .PAD(R_DATA[72]));
    INBUF \W_DATA_ibuf[42]  (.PAD(W_DATA[42]), .Y(W_DATA_c[42]));
    INBUF \W_DATA_ibuf[30]  (.PAD(W_DATA[30]), .Y(W_DATA_c[30]));
    OUTBUF \data_64_out_obuf[19]  (.D(W_DATA_c[23]), .PAD(
        data_64_out[19]));
    INBUF \selectt_ibuf[29]  (.PAD(selectt[29]), .Y(selectt_c[29]));
    error_gen error_gen_0 (.data_64_out_net_0({data_64_out_net_0[63], 
        data_64_out_net_0[62], data_64_out_net_0[61], 
        data_64_out_net_0[60], data_64_out_net_0[59], 
        data_64_out_net_0[58], data_64_out_net_0[57], 
        data_64_out_net_0[56], data_64_out_net_0[55], 
        data_64_out_net_0[54], data_64_out_net_0[53], 
        data_64_out_net_0[52], data_64_out_net_0[51], 
        data_64_out_net_0[50], data_64_out_net_0[49], 
        data_64_out_net_0[48], data_64_out_net_0[47], 
        data_64_out_net_0[46], data_64_out_net_0[45], 
        data_64_out_net_0[44], data_64_out_net_0[43], 
        data_64_out_net_0[42], data_64_out_net_0[41], 
        data_64_out_net_0[40], data_64_out_net_0[39], 
        data_64_out_net_0[38], data_64_out_net_0[37], 
        data_64_out_net_0[36], data_64_out_net_0[35], 
        data_64_out_net_0[34], data_64_out_net_0[33], 
        data_64_out_net_0[32], data_64_out_net_0[31], 
        data_64_out_net_0[30], data_64_out_net_0[29], 
        data_64_out_net_0[28], data_64_out_net_0[27], 
        data_64_out_net_0[26], data_64_out_net_0[25], 
        data_64_out_net_0[24], data_64_out_net_0[23], 
        data_64_out_net_0[22], data_64_out_net_0[21], 
        data_64_out_net_0[20], data_64_out_net_0[19], 
        data_64_out_net_0[18], data_64_out_net_0[17], 
        data_64_out_net_0[16], data_64_out_net_0[15], 
        data_64_out_net_0[14], data_64_out_net_0[13], 
        data_64_out_net_0[12], data_64_out_net_0[11], 
        data_64_out_net_0[10], data_64_out_net_0[9], 
        data_64_out_net_0[8], data_64_out_net_0[7], 
        data_64_out_net_0[6], data_64_out_net_0[5], 
        data_64_out_net_0[4], data_64_out_net_0[3], 
        data_64_out_net_0[2], data_64_out_net_0[1], 
        data_64_out_net_0[0]}), .R_DATA_c({R_DATA_c[77], R_DATA_c[76], 
        R_DATA_c[75], R_DATA_c[74], R_DATA_c[73], R_DATA_c[72], 
        R_DATA_c[71], R_DATA_c[70], N_51, N_50, R_DATA_c[67], 
        R_DATA_c[66], R_DATA_c[65], R_DATA_c[64], R_DATA_c[63], 
        R_DATA_c[62], R_DATA_c[61], R_DATA_c[60], N_49, N_48, 
        R_DATA_c[57], R_DATA_c[56], R_DATA_c[55], R_DATA_c[54], 
        R_DATA_c[53], R_DATA_c[52], R_DATA_c[51], R_DATA_c[50], N_47, 
        N_46, R_DATA_c[47], R_DATA_c[46], R_DATA_c[45], R_DATA_c[44], 
        R_DATA_c[43], R_DATA_c[42], R_DATA_c[41], R_DATA_c[40], N_45, 
        N_44, R_DATA_c[37], R_DATA_c[36], R_DATA_c[35], R_DATA_c[34], 
        R_DATA_c[33], R_DATA_c[32], R_DATA_c[31], R_DATA_c[30], N_43, 
        N_42, R_DATA_c[27], R_DATA_c[26], R_DATA_c[25], R_DATA_c[24], 
        R_DATA_c[23], R_DATA_c[22], R_DATA_c[21], R_DATA_c[20], N_41, 
        N_40, R_DATA_c[17], R_DATA_c[16], R_DATA_c[15], R_DATA_c[14], 
        R_DATA_c[13], R_DATA_c[12], R_DATA_c[11], R_DATA_c[10], N_39, 
        N_38, R_DATA_c[7], R_DATA_c[6], R_DATA_c[5], R_DATA_c[4], 
        R_DATA_c[3], R_DATA_c[2], R_DATA_c[1], R_DATA_c[0]}), 
        .selectt_c({selectt_c[63], selectt_c[62], selectt_c[61], 
        selectt_c[60], selectt_c[59], selectt_c[58], selectt_c[57], 
        selectt_c[56], selectt_c[55], selectt_c[54], selectt_c[53], 
        selectt_c[52], selectt_c[51], selectt_c[50], selectt_c[49], 
        selectt_c[48], selectt_c[47], selectt_c[46], selectt_c[45], 
        selectt_c[44], selectt_c[43], selectt_c[42], selectt_c[41], 
        selectt_c[40], selectt_c[39], selectt_c[38], selectt_c[37], 
        selectt_c[36], selectt_c[35], selectt_c[34], selectt_c[33], 
        selectt_c[32], selectt_c[31], selectt_c[30], selectt_c[29], 
        selectt_c[28], selectt_c[27], selectt_c[26], selectt_c[25], 
        selectt_c[24], selectt_c[23], selectt_c[22], selectt_c[21], 
        selectt_c[20], selectt_c[19], selectt_c[18], selectt_c[17], 
        selectt_c[16], selectt_c[15], selectt_c[14], selectt_c[13], 
        selectt_c[12], selectt_c[11], selectt_c[10], selectt_c[9], 
        selectt_c[8], selectt_c[7], selectt_c[6], selectt_c[5], 
        selectt_c[4], selectt_c[3], selectt_c[2], selectt_c[1], 
        selectt_c[0]}));
    OUTBUF \error_data_obuf[30]  (.D(error_data_c[30]), .PAD(
        error_data[30]));
    OUTBUF \data_64_out_obuf[49]  (.D(W_DATA_c[61]), .PAD(
        data_64_out[49]));
    OUTBUF \R_DATA_obuf[39]  (.D(R_DATA_c[39]), .PAD(R_DATA[39]));
    OUTBUF \R_DATA_obuf[1]  (.D(R_DATA_c[1]), .PAD(R_DATA[1]));
    INBUF \W_ADDR_ibuf[9]  (.PAD(W_ADDR[9]), .Y(W_ADDR_c[9]));
    OUTBUF \error_address_obuf[3]  (.D(error_address_c[3]), .PAD(
        error_address[3]));
    INBUF \W_ADDR_ibuf[13]  (.PAD(W_ADDR[13]), .Y(W_ADDR_c[13]));
    INBUF \W_DATA_ibuf[48]  (.PAD(W_DATA[48]), .Y(W_DATA_c[48]));
    OUTBUF \R_DATA_obuf[57]  (.D(R_DATA_c[57]), .PAD(R_DATA[57]));
    INBUF \R_ADDR_ibuf[3]  (.PAD(R_ADDR[3]), .Y(R_ADDR_c[3]));
    OUTBUF \R_DATA_obuf[36]  (.D(R_DATA_c[36]), .PAD(R_DATA[36]));
    INBUF \W_DATA_ibuf[46]  (.PAD(W_DATA[46]), .Y(W_DATA_c[46]));
    INBUF \selectt_ibuf[28]  (.PAD(selectt[28]), .Y(selectt_c[28]));
    INBUF \selectt_ibuf[20]  (.PAD(selectt[20]), .Y(selectt_c[20]));
    INBUF \WBYTE_EN_ibuf[0]  (.PAD(WBYTE_EN[0]), .Y(WBYTE_EN_c[0]));
    OUTBUF \error_data_obuf[55]  (.D(error_data_c[55]), .PAD(
        error_data[55]));
    OUTBUF \R_DATA_obuf[50]  (.D(R_DATA_c[50]), .PAD(R_DATA[50]));
    OUTBUF \error_data_obuf[33]  (.D(error_data_c[33]), .PAD(
        error_data[33]));
    OUTBUF \error_data_obuf[11]  (.D(error_data_c[11]), .PAD(
        error_data[11]));
    INBUF \W_DATA_ibuf[79]  (.PAD(W_DATA[79]), .Y(W_DATA_c[79]));
    OUTBUF \error_data_obuf[54]  (.D(error_data_c[54]), .PAD(
        error_data[54]));
    INBUF \W_DATA_ibuf[61]  (.PAD(W_DATA[61]), .Y(W_DATA_c[61]));
    INBUF \W_DATA_ibuf[5]  (.PAD(W_DATA[5]), .Y(W_DATA_c[5]));
    OUTBUF \data_64_out_obuf[52]  (.D(W_DATA_c[64]), .PAD(
        data_64_out[52]));
    INBUF \selectt_ibuf[24]  (.PAD(selectt[24]), .Y(selectt_c[24]));
    OUTBUF \R_DATA_obuf[69]  (.D(R_DATA_c[69]), .PAD(R_DATA[69]));
    OUTBUF \data_64_out_obuf[23]  (.D(W_DATA_c[27]), .PAD(
        data_64_out[23]));
    OUTBUF \error_address_obuf[13]  (.D(error_address_c[13]), .PAD(
        error_address[13]));
    INBUF \selectt_ibuf[42]  (.PAD(selectt[42]), .Y(selectt_c[42]));
    OUTBUF \error_data_obuf[9]  (.D(error_data_c[9]), .PAD(
        error_data[9]));
    INBUF \selectt_ibuf[47]  (.PAD(selectt[47]), .Y(selectt_c[47]));
    INBUF \selectt_ibuf[46]  (.PAD(selectt[46]), .Y(selectt_c[46]));
    INBUF \selectt_ibuf[63]  (.PAD(selectt[63]), .Y(selectt_c[63]));
    INBUF \W_DATA_ibuf[0]  (.PAD(W_DATA[0]), .Y(W_DATA_c[0]));
    OUTBUF \R_DATA_obuf[66]  (.D(R_DATA_c[66]), .PAD(R_DATA[66]));
    INBUF \R_ADDR_ibuf[5]  (.PAD(R_ADDR[5]), .Y(R_ADDR_c[5]));
    OUTBUF \error_data_obuf[47]  (.D(error_data_c[47]), .PAD(
        error_data[47]));
    OUTBUF \error_data_obuf[39]  (.D(error_data_c[39]), .PAD(
        error_data[39]));
    OUTBUF \data_64_out_obuf[30]  (.D(W_DATA_c[36]), .PAD(
        data_64_out[30]));
    OUTBUF \data_64_out_obuf[12]  (.D(W_DATA_c[14]), .PAD(
        data_64_out[12]));
    INBUF \W_DATA_ibuf[77]  (.PAD(W_DATA[77]), .Y(W_DATA_c[77]));
    OUTBUF \R_DATA_obuf[52]  (.D(R_DATA_c[52]), .PAD(R_DATA[52]));
    INBUF \W_DATA_ibuf[41]  (.PAD(W_DATA[41]), .Y(W_DATA_c[41]));
    OUTBUF \data_64_out_obuf[42]  (.D(W_DATA_c[52]), .PAD(
        data_64_out[42]));
    INBUF \selectt_ibuf[53]  (.PAD(selectt[53]), .Y(selectt_c[53]));
    OUTBUF \R_DATA_obuf[7]  (.D(R_DATA_c[7]), .PAD(R_DATA[7]));
    OUTBUF \R_DATA_obuf[75]  (.D(R_DATA_c[75]), .PAD(R_DATA[75]));
    OUTBUF \error_data_obuf[61]  (.D(error_data_c[61]), .PAD(
        error_data[61]));
    OUTBUF \data_64_out_obuf[9]  (.D(W_DATA_c[11]), .PAD(
        data_64_out[9]));
    OUTBUF error_flag_obuf (.D(ERRr_c), .PAD(error_flag));
    OUTBUF \error_address_obuf[12]  (.D(error_address_c[12]), .PAD(
        error_address[12]));
    INBUF \selectt_ibuf[15]  (.PAD(selectt[15]), .Y(selectt_c[15]));
    OUTBUF \data_64_out_obuf[63]  (.D(W_DATA_c[77]), .PAD(
        data_64_out[63]));
    INBUF \W_DATA_ibuf[29]  (.PAD(W_DATA[29]), .Y(W_DATA_c[29]));
    INBUF \R_ADDR_ibuf[12]  (.PAD(R_ADDR[12]), .Y(R_ADDR_c[12]));
    OUTBUF \error_data_obuf[16]  (.D(error_data_c[16]), .PAD(
        error_data[16]));
    INBUF \W_DATA_ibuf[59]  (.PAD(W_DATA[59]), .Y(W_DATA_c[59]));
    OUTBUF \error_data_obuf[51]  (.D(error_data_c[51]), .PAD(
        error_data[51]));
    OUTBUF \R_DATA_obuf[73]  (.D(R_DATA_c[73]), .PAD(R_DATA[73]));
    INBUF \W_DATA_ibuf[63]  (.PAD(W_DATA[63]), .Y(W_DATA_c[63]));
    INBUF \W_ADDR_ibuf[0]  (.PAD(W_ADDR[0]), .Y(W_ADDR_c[0]));
    OUTBUF \error_data_obuf[12]  (.D(error_data_c[12]), .PAD(
        error_data[12]));
    OUTBUF \data_64_out_obuf[29]  (.D(W_DATA_c[35]), .PAD(
        data_64_out[29]));
    INBUF \W_DATA_ibuf[8]  (.PAD(W_DATA[8]), .Y(W_DATA_c[8]));
    OUTBUF \data_64_out_obuf[31]  (.D(W_DATA_c[37]), .PAD(
        data_64_out[31]));
    OUTBUF \R_DATA_obuf[3]  (.D(R_DATA_c[3]), .PAD(R_DATA[3]));
    INBUF \W_DATA_ibuf[3]  (.PAD(W_DATA[3]), .Y(W_DATA_c[3]));
    INBUF \W_DATA_ibuf[27]  (.PAD(W_DATA[27]), .Y(W_DATA_c[27]));
    OUTBUF \R_DATA_obuf[74]  (.D(R_DATA_c[74]), .PAD(R_DATA[74]));
    INBUF \W_DATA_ibuf[57]  (.PAD(W_DATA[57]), .Y(W_DATA_c[57]));
    INBUF R_EN_ibuf (.PAD(R_EN), .Y(R_EN_c));
    INBUF \WBYTE_EN_ibuf[2]  (.PAD(WBYTE_EN[2]), .Y(WBYTE_EN_c[2]));
    INBUF \selectt_ibuf[21]  (.PAD(selectt[21]), .Y(selectt_c[21]));
    OUTBUF \error_data_obuf[40]  (.D(error_data_c[40]), .PAD(
        error_data[40]));
    INBUF \W_DATA_ibuf[43]  (.PAD(W_DATA[43]), .Y(W_DATA_c[43]));
    OUTBUF \error_data_obuf[28]  (.D(error_data_c[28]), .PAD(
        error_data[28]));
    INBUF \W_ADDR_ibuf[1]  (.PAD(W_ADDR[1]), .Y(W_ADDR_c[1]));
    INBUF \selectt_ibuf[49]  (.PAD(selectt[49]), .Y(selectt_c[49]));
    INBUF \W_DATA_ibuf[19]  (.PAD(W_DATA[19]), .Y(W_DATA_c[19]));
    CLKINT I_1 (.A(CLK_ibuf_Z), .Y(NN_1));
    OUTBUF \R_DATA_obuf[78]  (.D(R_DATA_c[78]), .PAD(R_DATA[78]));
    OUTBUF \data_64_out_obuf[54]  (.D(W_DATA_c[66]), .PAD(
        data_64_out[54]));
    INBUF \R_ADDR_ibuf[2]  (.PAD(R_ADDR[2]), .Y(R_ADDR_c[2]));
    OUTBUF \error_data_obuf[62]  (.D(error_data_c[62]), .PAD(
        error_data[62]));
    OUTBUF \error_address_obuf[5]  (.D(error_address_c[5]), .PAD(
        error_address[5]));
    OUTBUF \R_DATA_obuf[47]  (.D(R_DATA_c[47]), .PAD(R_DATA[47]));
    INBUF \W_DATA_ibuf[39]  (.PAD(W_DATA[39]), .Y(W_DATA_c[39]));
    OUTBUF \error_data_obuf[35]  (.D(error_data_c[35]), .PAD(
        error_data[35]));
    OUTBUF \R_DATA_obuf[9]  (.D(R_DATA_c[9]), .PAD(R_DATA[9]));
    OUTBUF \R_DATA_obuf[8]  (.D(R_DATA_c[8]), .PAD(R_DATA[8]));
    OUTBUF \error_data_obuf[56]  (.D(error_data_c[56]), .PAD(
        error_data[56]));
    OUTBUF \error_data_obuf[43]  (.D(error_data_c[43]), .PAD(
        error_data[43]));
    OUTBUF \R_DATA_obuf[71]  (.D(R_DATA_c[71]), .PAD(R_DATA[71]));
    INBUF \selectt_ibuf[48]  (.PAD(selectt[48]), .Y(selectt_c[48]));
    OUTBUF \R_DATA_obuf[55]  (.D(R_DATA_c[55]), .PAD(R_DATA[55]));
    OUTBUF \R_DATA_obuf[40]  (.D(R_DATA_c[40]), .PAD(R_DATA[40]));
    OUTBUF \error_data_obuf[52]  (.D(error_data_c[52]), .PAD(
        error_data[52]));
    OUTBUF \error_data_obuf[34]  (.D(error_data_c[34]), .PAD(
        error_data[34]));
    INBUF \selectt_ibuf[40]  (.PAD(selectt[40]), .Y(selectt_c[40]));
    INBUF \W_DATA_ibuf[17]  (.PAD(W_DATA[17]), .Y(W_DATA_c[17]));
    INBUF \W_DATA_ibuf[72]  (.PAD(W_DATA[72]), .Y(W_DATA_c[72]));
    INBUF \W_DATA_ibuf[9]  (.PAD(W_DATA[9]), .Y(W_DATA_c[9]));
    OUTBUF \data_64_out_obuf[38]  (.D(W_DATA_c[46]), .PAD(
        data_64_out[38]));
    OUTBUF \data_64_out_obuf[14]  (.D(W_DATA_c[16]), .PAD(
        data_64_out[14]));
    INBUF \selectt_ibuf[7]  (.PAD(selectt[7]), .Y(selectt_c[7]));
    INBUF \selectt_ibuf[12]  (.PAD(selectt[12]), .Y(selectt_c[12]));
    INBUF \selectt_ibuf[17]  (.PAD(selectt[17]), .Y(selectt_c[17]));
    INBUF \selectt_ibuf[16]  (.PAD(selectt[16]), .Y(selectt_c[16]));
    OUTBUF \data_64_out_obuf[22]  (.D(W_DATA_c[26]), .PAD(
        data_64_out[22]));
    INBUF \W_DATA_ibuf[37]  (.PAD(W_DATA[37]), .Y(W_DATA_c[37]));
    OUTBUF \R_DATA_obuf[53]  (.D(R_DATA_c[53]), .PAD(R_DATA[53]));
    INBUF \WBYTE_EN_ibuf[1]  (.PAD(WBYTE_EN[1]), .Y(WBYTE_EN_c[1]));
    INBUF \selectt_ibuf[9]  (.PAD(selectt[9]), .Y(selectt_c[9]));
    OUTBUF \data_64_out_obuf[44]  (.D(W_DATA_c[54]), .PAD(
        data_64_out[44]));
    INBUF \selectt_ibuf[44]  (.PAD(selectt[44]), .Y(selectt_c[44]));
    INBUF \selectt_ibuf[35]  (.PAD(selectt[35]), .Y(selectt_c[35]));
    OUTBUF \error_data_obuf[4]  (.D(error_data_c[4]), .PAD(
        error_data[4]));
    INBUF \W_ADDR_ibuf[11]  (.PAD(W_ADDR[11]), .Y(W_ADDR_c[11]));
    PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM 
        PF_SRAM_AHBL_AXI_C1_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_0 (.R_DATA_c({
        R_DATA_c[79], R_DATA_c[78], R_DATA_c[77], R_DATA_c[76], 
        R_DATA_c[75], R_DATA_c[74], R_DATA_c[73], R_DATA_c[72], 
        R_DATA_c[71], R_DATA_c[70], R_DATA_c[69], R_DATA_c[68], 
        R_DATA_c[67], R_DATA_c[66], R_DATA_c[65], R_DATA_c[64], 
        R_DATA_c[63], R_DATA_c[62], R_DATA_c[61], R_DATA_c[60], 
        R_DATA_c[59], R_DATA_c[58], R_DATA_c[57], R_DATA_c[56], 
        R_DATA_c[55], R_DATA_c[54], R_DATA_c[53], R_DATA_c[52], 
        R_DATA_c[51], R_DATA_c[50], R_DATA_c[49], R_DATA_c[48], 
        R_DATA_c[47], R_DATA_c[46], R_DATA_c[45], R_DATA_c[44], 
        R_DATA_c[43], R_DATA_c[42], R_DATA_c[41], R_DATA_c[40], 
        R_DATA_c[39], R_DATA_c[38], R_DATA_c[37], R_DATA_c[36], 
        R_DATA_c[35], R_DATA_c[34], R_DATA_c[33], R_DATA_c[32], 
        R_DATA_c[31], R_DATA_c[30], R_DATA_c[29], R_DATA_c[28], 
        R_DATA_c[27], R_DATA_c[26], R_DATA_c[25], R_DATA_c[24], 
        R_DATA_c[23], R_DATA_c[22], R_DATA_c[21], R_DATA_c[20], 
        R_DATA_c[19], R_DATA_c[18], R_DATA_c[17], R_DATA_c[16], 
        R_DATA_c[15], R_DATA_c[14], R_DATA_c[13], R_DATA_c[12], 
        R_DATA_c[11], R_DATA_c[10], R_DATA_c[9], R_DATA_c[8], 
        R_DATA_c[7], R_DATA_c[6], R_DATA_c[5], R_DATA_c[4], 
        R_DATA_c[3], R_DATA_c[2], R_DATA_c[1], R_DATA_c[0]}), 
        .WBYTE_EN_c({WBYTE_EN_c[7], WBYTE_EN_c[6], WBYTE_EN_c[5], 
        WBYTE_EN_c[4], WBYTE_EN_c[3], WBYTE_EN_c[2], WBYTE_EN_c[1], 
        WBYTE_EN_c[0]}), .W_DATA_c({W_DATA_c[79], W_DATA_c[78], 
        W_DATA_c[77], W_DATA_c[76], W_DATA_c[75], W_DATA_c[74], 
        W_DATA_c[73], W_DATA_c[72], W_DATA_c[71], W_DATA_c[70], 
        W_DATA_c[69], W_DATA_c[68], W_DATA_c[67], W_DATA_c[66], 
        W_DATA_c[65], W_DATA_c[64], W_DATA_c[63], W_DATA_c[62], 
        W_DATA_c[61], W_DATA_c[60], W_DATA_c[59], W_DATA_c[58], 
        W_DATA_c[57], W_DATA_c[56], W_DATA_c[55], W_DATA_c[54], 
        W_DATA_c[53], W_DATA_c[52], W_DATA_c[51], W_DATA_c[50], 
        W_DATA_c[49], W_DATA_c[48], W_DATA_c[47], W_DATA_c[46], 
        W_DATA_c[45], W_DATA_c[44], W_DATA_c[43], W_DATA_c[42], 
        W_DATA_c[41], W_DATA_c[40], W_DATA_c[39], W_DATA_c[38], 
        W_DATA_c[37], W_DATA_c[36], W_DATA_c[35], W_DATA_c[34], 
        W_DATA_c[33], W_DATA_c[32], W_DATA_c[31], W_DATA_c[30], 
        W_DATA_c[29], W_DATA_c[28], W_DATA_c[27], W_DATA_c[26], 
        W_DATA_c[25], W_DATA_c[24], W_DATA_c[23], W_DATA_c[22], 
        W_DATA_c[21], W_DATA_c[20], W_DATA_c[19], W_DATA_c[18], 
        W_DATA_c[17], W_DATA_c[16], W_DATA_c[15], W_DATA_c[14], 
        W_DATA_c[13], W_DATA_c[12], W_DATA_c[11], W_DATA_c[10], 
        W_DATA_c[9], W_DATA_c[8], W_DATA_c[7], W_DATA_c[6], 
        W_DATA_c[5], W_DATA_c[4], W_DATA_c[3], W_DATA_c[2], 
        W_DATA_c[1], W_DATA_c[0]}), .W_ADDR_c({W_ADDR_c[13], 
        W_ADDR_c[12], W_ADDR_c[11], W_ADDR_c[10], W_ADDR_c[9], 
        W_ADDR_c[8], W_ADDR_c[7], W_ADDR_c[6], W_ADDR_c[5], 
        W_ADDR_c[4], W_ADDR_c[3], W_ADDR_c[2], W_ADDR_c[1], 
        W_ADDR_c[0]}), .R_ADDR_c({R_ADDR_c[13], R_ADDR_c[12], 
        R_ADDR_c[11], R_ADDR_c[10], R_ADDR_c[9], R_ADDR_c[8], 
        R_ADDR_c[7], R_ADDR_c[6], R_ADDR_c[5], R_ADDR_c[4], 
        R_ADDR_c[3], R_ADDR_c[2], R_ADDR_c[1], R_ADDR_c[0]}), .CLK(
        NN_1), .R_EN_c(R_EN_c), .W_EN_c(W_EN_c));
    OUTBUF \error_data_obuf[49]  (.D(error_data_c[49]), .PAD(
        error_data[49]));
    INBUF \W_DATA_ibuf[78]  (.PAD(W_DATA[78]), .Y(W_DATA_c[78]));
    OUTBUF \R_DATA_obuf[17]  (.D(R_DATA_c[17]), .PAD(R_DATA[17]));
    INBUF \R_ADDR_ibuf[8]  (.PAD(R_ADDR[8]), .Y(R_ADDR_c[8]));
    INBUF \W_DATA_ibuf[64]  (.PAD(W_DATA[64]), .Y(W_DATA_c[64]));
    OUTBUF \R_DATA_obuf[27]  (.D(R_DATA_c[27]), .PAD(R_DATA[27]));
    INBUF \W_DATA_ibuf[76]  (.PAD(W_DATA[76]), .Y(W_DATA_c[76]));
    OUTBUF \R_DATA_obuf[54]  (.D(R_DATA_c[54]), .PAD(R_DATA[54]));
    OUTBUF \error_data_obuf[0]  (.D(error_data_c[0]), .PAD(
        error_data[0]));
    OUTBUF \R_DATA_obuf[42]  (.D(R_DATA_c[42]), .PAD(R_DATA[42]));
    OUTBUF \error_data_obuf[8]  (.D(error_data_c[8]), .PAD(
        error_data[8]));
    OUTBUF \R_DATA_obuf[10]  (.D(R_DATA_c[10]), .PAD(R_DATA[10]));
    OUTBUF \R_DATA_obuf[5]  (.D(R_DATA_c[5]), .PAD(R_DATA[5]));
    OUTBUF \R_DATA_obuf[20]  (.D(R_DATA_c[20]), .PAD(R_DATA[20]));
    INBUF \R_ADDR_ibuf[0]  (.PAD(R_ADDR[0]), .Y(R_ADDR_c[0]));
    OUTBUF \R_DATA_obuf[0]  (.D(R_DATA_c[0]), .PAD(R_DATA[0]));
    OUTBUF \error_data_obuf[31]  (.D(error_data_c[31]), .PAD(
        error_data[31]));
    OUTBUF \data_64_out_obuf[62]  (.D(W_DATA_c[76]), .PAD(
        data_64_out[62]));
    INBUF \W_DATA_ibuf[22]  (.PAD(W_DATA[22]), .Y(W_DATA_c[22]));
    OUTBUF \error_data_obuf[27]  (.D(error_data_c[27]), .PAD(
        error_data[27]));
    INBUF \W_DATA_ibuf[52]  (.PAD(W_DATA[52]), .Y(W_DATA_c[52]));
    OUTBUF \R_DATA_obuf[58]  (.D(R_DATA_c[58]), .PAD(R_DATA[58]));
    INBUF \W_DATA_ibuf[44]  (.PAD(W_DATA[44]), .Y(W_DATA_c[44]));
    INBUF \selectt_ibuf[23]  (.PAD(selectt[23]), .Y(selectt_c[23]));
    OUTBUF \data_64_out_obuf[50]  (.D(W_DATA_c[62]), .PAD(
        data_64_out[50]));
    OUTBUF \R_DATA_obuf[51]  (.D(R_DATA_c[51]), .PAD(R_DATA[51]));
    INBUF \W_ADDR_ibuf[4]  (.PAD(W_ADDR[4]), .Y(W_ADDR_c[4]));
    INBUF \selectt_ibuf[8]  (.PAD(selectt[8]), .Y(selectt_c[8]));
    INBUF \W_DATA_ibuf[28]  (.PAD(W_DATA[28]), .Y(W_DATA_c[28]));
    OUTBUF \R_DATA_obuf[12]  (.D(R_DATA_c[12]), .PAD(R_DATA[12]));
    OUTBUF \R_DATA_obuf[79]  (.D(R_DATA_c[79]), .PAD(R_DATA[79]));
    OUTBUF \R_DATA_obuf[22]  (.D(R_DATA_c[22]), .PAD(R_DATA[22]));
    INBUF \W_DATA_ibuf[71]  (.PAD(W_DATA[71]), .Y(W_DATA_c[71]));
    INBUF \W_DATA_ibuf[58]  (.PAD(W_DATA[58]), .Y(W_DATA_c[58]));
    OUTBUF \data_64_out_obuf[10]  (.D(W_DATA_c[12]), .PAD(
        data_64_out[10]));
    INBUF \W_DATA_ibuf[26]  (.PAD(W_DATA[26]), .Y(W_DATA_c[26]));
    OUTBUF \error_data_obuf[5]  (.D(error_data_c[5]), .PAD(
        error_data[5]));
    INBUF \W_DATA_ibuf[56]  (.PAD(W_DATA[56]), .Y(W_DATA_c[56]));
    INBUF \selectt_ibuf[19]  (.PAD(selectt[19]), .Y(selectt_c[19]));
    INBUF \R_ADDR_ibuf[1]  (.PAD(R_ADDR[1]), .Y(R_ADDR_c[1]));
    OUTBUF \data_64_out_obuf[35]  (.D(W_DATA_c[43]), .PAD(
        data_64_out[35]));
    
endmodule
