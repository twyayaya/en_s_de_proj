///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: test1_tb.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::PolarFire> <Die::MPF300TS> <Package::FCG1152>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

`timescale 1ns/100ps

module test1_tb;

parameter SYSCLK_PERIOD = 100;// 10MHZ

reg SYSCLK;
reg NSYSRESET;

initial
begin
    SYSCLK = 1'b0;
    NSYSRESET = 1'b0;
end

//////////////////////////////////////////////////////////////////////
// Reset Pulse
//////////////////////////////////////////////////////////////////////
initial
begin
    #(SYSCLK_PERIOD * 10 )
        NSYSRESET = 1'b1;
end


//////////////////////////////////////////////////////////////////////
// Clock Driver
//////////////////////////////////////////////////////////////////////
always @(SYSCLK)
    #(SYSCLK_PERIOD / 2.0) SYSCLK <= !SYSCLK;


//////////////////////////////////////////////////////////////////////
// Instantiate Unit Under Test:  test1
//////////////////////////////////////////////////////////////////////

reg [71:0] INn;

wire [63:0] real_data;
wire ERRr;

test1 test1_0 (
    // Inputs
    .clk(SYSCLK),
    .INn(INn),

    // Outputs
    .real_data(real_data),
    .ERRr(ERRr)


);

initial begin
#50
INn = 72'b000000000000000000000000000000000000000000000000000000000000000000000001;//1
#10
INn = 72'b010110100001000111000110110000110101000100001101110000001000001000011010;//2
#10
INn = 72'b001001100010110110111011001100000110111100010000111001011111001110111011;//3
#10
INn = 72'b101100110110010000100110000100101011010000010111010000000011110010111001;//4
#10
INn = 72'b101111000100111001011100111110011111100111100000100000011000001110000110;//12
#10
INn = 72'b000011110100001100011001101111001010001001001111000000000101011010010001;//34
#10
INn = 72'b111100110101011111100011110111000000111001111001010011100000001000101110;
#10
INn = 72'b100100010110101010101001110100001101010010100000110001011100111001011101;
#10
INn = 72'b000001100011100000111010101111011011000100111001011101001111101111101011;
#10
INn = 72'b111001110110110100000100111110010000100110011101110110001100100000011000;


end


initial begin
    $monitor($time, ": real_data = %b, real_data = %d ,  ERRr = %b", real_data, real_data, ERRr  );
end

endmodule

