`timescale 1ns / 100ps


module error_gen_for_72bit(
    input [71:0] INn,
    output [71:0] OUTt,
    input [63:0] selectt
    );
    
reg [71:0] IN_2;



always@(*) begin
    IN_2 = INn;
    case(selectt)
        64'd0  : IN_2[0] = ~INn[0] ;
        64'd1  : IN_2[1] = ~INn[1] ;
        64'd2  : IN_2[2] = ~INn[2] ;
        64'd3  : IN_2[3] = ~INn[3] ;
        64'd4  : IN_2[4] = ~INn[4] ;
        64'd5  : IN_2[5] = ~INn[5] ;
        64'd6  : IN_2[6] = ~INn[6] ;
        64'd7  : IN_2[7] = ~INn[7] ;
        64'd8  : IN_2[8] = ~INn[8] ;
        64'd9  : IN_2[9] = ~INn[9] ;
        64'd10  : IN_2[10] = ~INn[10] ;
        64'd11  : IN_2[11] = ~INn[11] ;
        64'd12  : IN_2[12] = ~INn[12] ;
        64'd13  : IN_2[13] = ~INn[13] ;
        64'd14  : IN_2[14] = ~INn[14] ;
        64'd15  : IN_2[15] = ~INn[15] ;
        64'd16  : IN_2[16] = ~INn[16] ;
        64'd17  : IN_2[17] = ~INn[17] ;
        64'd18  : IN_2[18] = ~INn[18] ;
        64'd19  : IN_2[19] = ~INn[19] ;
        64'd20  : IN_2[20] = ~INn[20] ;
        64'd21  : IN_2[21] = ~INn[21] ;
        64'd22  : IN_2[22] = ~INn[22] ;
        64'd23  : IN_2[23] = ~INn[23] ;
        64'd24  : IN_2[24] = ~INn[24] ;
        64'd25  : IN_2[25] = ~INn[25] ;
        64'd26  : IN_2[26] = ~INn[26] ;
        64'd27  : IN_2[27] = ~INn[27] ;
        64'd28  : IN_2[28] = ~INn[28] ;
        64'd29  : IN_2[29] = ~INn[29] ;
        64'd30  : IN_2[30] = ~INn[30] ;
        64'd31  : IN_2[31] = ~INn[31] ;
        64'd32  : IN_2[32] = ~INn[32] ;
        64'd33  : IN_2[33] = ~INn[33] ;
        64'd34  : IN_2[34] = ~INn[34] ;
        64'd35  : IN_2[35] = ~INn[35] ;
        64'd36  : IN_2[36] = ~INn[36] ;
        64'd37  : IN_2[37] = ~INn[37] ;
        64'd38  : IN_2[38] = ~INn[38] ;
        64'd39  : IN_2[39] = ~INn[39] ;
        64'd40  : IN_2[40] = ~INn[40] ;
        64'd41  : IN_2[41] = ~INn[41] ;
        64'd42  : IN_2[42] = ~INn[42] ;
        64'd43  : IN_2[43] = ~INn[43] ;
        64'd44  : IN_2[44] = ~INn[44] ;
        64'd45  : IN_2[45] = ~INn[45] ;
        64'd46  : IN_2[46] = ~INn[46] ;
        64'd47  : IN_2[47] = ~INn[47] ;
        64'd48  : IN_2[48] = ~INn[48] ;
        64'd49  : IN_2[49] = ~INn[49] ;
        64'd50  : IN_2[50] = ~INn[50] ;
        64'd51  : IN_2[51] = ~INn[51] ;
        64'd52  : IN_2[52] = ~INn[52] ;
        64'd53  : IN_2[53] = ~INn[53] ;
        64'd54  : IN_2[54] = ~INn[54] ;
        64'd55  : IN_2[55] = ~INn[55] ;
        64'd56  : IN_2[56] = ~INn[56] ;
        64'd57  : IN_2[57] = ~INn[57] ;
        64'd58  : IN_2[58] = ~INn[58] ;
        64'd59  : IN_2[59] = ~INn[59] ;
        64'd60  : IN_2[60] = ~INn[60] ;
        64'd61  : IN_2[61] = ~INn[61] ;
        64'd62  : IN_2[62] = ~INn[62] ;
        64'd63  : IN_2[63] = ~INn[63] ;
        
        default: IN_2 = INn ;
    endcase
end

assign OUTt = IN_2;

endmodule